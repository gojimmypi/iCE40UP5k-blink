-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 6 2018 12:49:44

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    RGB2 : out std_logic;
    RGB1 : out std_logic;
    RGB0 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2111\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \ctrZ0Z_0\ : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal \ctrZ0Z_1\ : std_logic;
signal ctr_cry_0 : std_logic;
signal \ctrZ0Z_2\ : std_logic;
signal ctr_cry_1 : std_logic;
signal \ctrZ0Z_3\ : std_logic;
signal ctr_cry_2 : std_logic;
signal \ctrZ0Z_4\ : std_logic;
signal ctr_cry_3 : std_logic;
signal \ctrZ0Z_5\ : std_logic;
signal ctr_cry_4 : std_logic;
signal \ctrZ0Z_6\ : std_logic;
signal ctr_cry_5 : std_logic;
signal \ctrZ0Z_7\ : std_logic;
signal ctr_cry_6 : std_logic;
signal ctr_cry_7 : std_logic;
signal \ctrZ0Z_8\ : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal \ctrZ0Z_9\ : std_logic;
signal ctr_cry_8 : std_logic;
signal \ctrZ0Z_10\ : std_logic;
signal ctr_cry_9 : std_logic;
signal \ctrZ0Z_11\ : std_logic;
signal ctr_cry_10 : std_logic;
signal \ctrZ0Z_12\ : std_logic;
signal ctr_cry_11 : std_logic;
signal \ctrZ0Z_13\ : std_logic;
signal ctr_cry_12 : std_logic;
signal \ctrZ0Z_14\ : std_logic;
signal ctr_cry_13 : std_logic;
signal \ctrZ0Z_15\ : std_logic;
signal ctr_cry_14 : std_logic;
signal ctr_cry_15 : std_logic;
signal \ctrZ0Z_16\ : std_logic;
signal \bfn_1_27_0_\ : std_logic;
signal \ctrZ0Z_17\ : std_logic;
signal ctr_cry_16 : std_logic;
signal ctr_cry_17 : std_logic;
signal ctr_cry_18 : std_logic;
signal ctr_cry_19 : std_logic;
signal ctr_cry_20 : std_logic;
signal ctr_cry_21 : std_logic;
signal ctr_cry_22 : std_logic;
signal ctr_cry_23 : std_logic;
signal \bfn_1_28_0_\ : std_logic;
signal ctr_cry_24 : std_logic;
signal ctr_cry_25 : std_logic;
signal ctr_cry_26 : std_logic;
signal ctr_cry_27 : std_logic;
signal ctr_cry_28 : std_logic;
signal ctr_cry_29 : std_logic;
signal ctr_cry_30 : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal pwm_ctr_cry_0 : std_logic;
signal pwm_ctr_cry_1 : std_logic;
signal pwm_ctr_cry_2 : std_logic;
signal pwm_ctr_cry_3 : std_logic;
signal pwm_ctr_cry_4 : std_logic;
signal pwm_ctr_cry_5 : std_logic;
signal pwm_ctr_cry_6 : std_logic;
signal pwm_ctr_cry_7 : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal pwm_ctr_cry_8 : std_logic;
signal pwm_ctr_cry_9 : std_logic;
signal pwm_ctr_cry_10 : std_logic;
signal \N_88_cascade_\ : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal un34_r_val_0_cry_1 : std_logic;
signal un34_r_val_0_cry_2 : std_logic;
signal un34_r_val_0_cry_3 : std_logic;
signal un34_r_val_0_cry_4 : std_logic;
signal un34_r_val_0_cry_5 : std_logic;
signal un34_r_val_0_cry_6 : std_logic;
signal un34_r_val_0_cry_7 : std_logic;
signal un34_r_val_0_cry_8 : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal un34_r_val_0_cry_9 : std_logic;
signal un34_r_val_0_cry_10 : std_logic;
signal \un34_r_val_0_cry_10_THRU_CO_cascade_\ : std_logic;
signal \N_92_cascade_\ : std_logic;
signal \N_66_cascade_\ : std_logic;
signal \N_87_cascade_\ : std_logic;
signal \ctrZ0Z_19\ : std_logic;
signal \un40_b_val_3_ns_1_1_cascade_\ : std_logic;
signal pwm_g_1_0 : std_logic;
signal \pwm_ctrZ0Z_0\ : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal \pwm_ctrZ0Z_1\ : std_logic;
signal pwm_g_1_1 : std_logic;
signal pwm_g_1_cry_0 : std_logic;
signal \pwm_ctrZ0Z_2\ : std_logic;
signal pwm_g_1_2 : std_logic;
signal pwm_g_1_cry_1 : std_logic;
signal \pwm_ctrZ0Z_3\ : std_logic;
signal pwm_g_1_3 : std_logic;
signal pwm_g_1_cry_2 : std_logic;
signal \pwm_ctrZ0Z_4\ : std_logic;
signal pwm_g_1_cry_3 : std_logic;
signal pwm_g_1_5 : std_logic;
signal \pwm_ctrZ0Z_5\ : std_logic;
signal pwm_g_1_cry_4 : std_logic;
signal \pwm_ctrZ0Z_6\ : std_logic;
signal pwm_g_1_cry_5 : std_logic;
signal \pwm_ctrZ0Z_7\ : std_logic;
signal pwm_g_1_cry_6 : std_logic;
signal pwm_g_1_cry_7 : std_logic;
signal pwm_g_1_8 : std_logic;
signal \pwm_ctrZ0Z_8\ : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal pwm_g_1_9 : std_logic;
signal \pwm_ctrZ0Z_9\ : std_logic;
signal pwm_g_1_cry_8 : std_logic;
signal \pwm_ctrZ0Z_10\ : std_logic;
signal pwm_g_1_cry_9 : std_logic;
signal \pwm_ctrZ0Z_11\ : std_logic;
signal pwm_g_1_11 : std_logic;
signal pwm_g_1_cry_10 : std_logic;
signal pwm_g_1 : std_logic;
signal \pwm_gZ0\ : std_logic;
signal \N_71_cascade_\ : std_logic;
signal pwm_g_1_10 : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \ctr_RNI7D9MZ0Z_21\ : std_logic;
signal \un33_r_val_cry_0_THRU_CO\ : std_logic;
signal un33_r_val_cry_0 : std_logic;
signal un33_r_val_cry_1 : std_logic;
signal un33_r_val_cry_2 : std_logic;
signal un33_r_val_cry_3 : std_logic;
signal \un33_r_val_cry_4_THRU_CO\ : std_logic;
signal un33_r_val_cry_4 : std_logic;
signal un33_r_val_cry_5 : std_logic;
signal un33_r_val_cry_6 : std_logic;
signal un33_r_val_cry_7 : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal un33_r_val_cry_8 : std_logic;
signal un33_r_val_cry_9 : std_logic;
signal un33_r_val_cry_10 : std_logic;
signal \un33_r_val_cry_10_THRU_CO_cascade_\ : std_logic;
signal \un34_r_val_0_cry_10_THRU_CO\ : std_logic;
signal \un33_r_val_cry_3_THRU_CO\ : std_logic;
signal \N_91_cascade_\ : std_logic;
signal pwm_r_1_0 : std_logic;
signal \bfn_3_27_0_\ : std_logic;
signal pwm_r_1_1 : std_logic;
signal pwm_r_1_cry_0 : std_logic;
signal pwm_r_1_cry_1 : std_logic;
signal pwm_r_1_cry_2 : std_logic;
signal pwm_r_1_4 : std_logic;
signal pwm_r_1_cry_3 : std_logic;
signal pwm_r_1_5 : std_logic;
signal pwm_r_1_cry_4 : std_logic;
signal pwm_r_1_cry_5 : std_logic;
signal pwm_r_1_cry_6 : std_logic;
signal pwm_r_1_cry_7 : std_logic;
signal \bfn_3_28_0_\ : std_logic;
signal pwm_r_1_cry_8 : std_logic;
signal pwm_r_1_cry_9 : std_logic;
signal pwm_r_1_cry_10 : std_logic;
signal pwm_r_1 : std_logic;
signal \pwm_rZ0\ : std_logic;
signal \un33_r_val_cry_8_THRU_CO\ : std_logic;
signal \N_96_cascade_\ : std_logic;
signal pwm_r_1_9 : std_logic;
signal \un34_r_val_0_cry_9_c_RNIV0HKZ0\ : std_logic;
signal pwm_ctr_i_0 : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal pwm_ctr_i_1 : std_logic;
signal pwm_b_1_1 : std_logic;
signal pwm_b_1_cry_0 : std_logic;
signal pwm_ctr_i_2 : std_logic;
signal pwm_b_1_cry_1 : std_logic;
signal pwm_b_1_3 : std_logic;
signal pwm_ctr_i_3 : std_logic;
signal pwm_b_1_cry_2 : std_logic;
signal pwm_ctr_i_4 : std_logic;
signal pwm_b_1_cry_3 : std_logic;
signal pwm_ctr_i_5 : std_logic;
signal pwm_b_1_cry_4 : std_logic;
signal pwm_ctr_i_6 : std_logic;
signal pwm_b_1_cry_5 : std_logic;
signal pwm_ctr_i_7 : std_logic;
signal pwm_b_1_cry_6 : std_logic;
signal pwm_b_1_cry_7 : std_logic;
signal pwm_b_1_8 : std_logic;
signal pwm_ctr_i_8 : std_logic;
signal \bfn_3_30_0_\ : std_logic;
signal pwm_ctr_i_9 : std_logic;
signal pwm_b_1_cry_8 : std_logic;
signal pwm_b_1_10 : std_logic;
signal pwm_ctr_i_10 : std_logic;
signal pwm_b_1_cry_9 : std_logic;
signal pwm_b_1_11 : std_logic;
signal pwm_ctr_i_11 : std_logic;
signal pwm_b_1_cry_10 : std_logic;
signal pwm_b_1 : std_logic;
signal \pwm_bZ0\ : std_logic;
signal clk : std_logic;
signal \un34_r_val_0_cry_8_c_RNI9TKVZ0\ : std_logic;
signal \N_72_cascade_\ : std_logic;
signal pwm_b_1_9 : std_logic;
signal \un33_r_val_cry_1_THRU_CO\ : std_logic;
signal \N_89_cascade_\ : std_logic;
signal pwm_r_1_2 : std_logic;
signal \ctrZ0Z_21\ : std_logic;
signal \un34_r_val_0_cry_2_c_RNIN4EVZ0\ : std_logic;
signal \un33_r_val_cry_2_THRU_CO\ : std_logic;
signal \N_90_cascade_\ : std_logic;
signal pwm_r_1_3 : std_logic;
signal \un33_r_val_cry_5_THRU_CO\ : std_logic;
signal \N_93_cascade_\ : std_logic;
signal pwm_r_1_6 : std_logic;
signal \ctrZ0Z_23\ : std_logic;
signal \un34_r_val_0_cry_4_c_RNITCGVZ0\ : std_logic;
signal \N_68_cascade_\ : std_logic;
signal pwm_b_1_5 : std_logic;
signal \un33_r_val_cry_6_THRU_CO\ : std_logic;
signal \N_94_cascade_\ : std_logic;
signal pwm_r_1_7 : std_logic;
signal \ctrZ0Z_29\ : std_logic;
signal \pwm_r_1_cry_11_c_RNOZ0Z_0\ : std_logic;
signal pwm_r_1_11 : std_logic;
signal pwm_g_1_6 : std_logic;
signal \un34_r_val_0_cry_7_c_RNI6PJVZ0\ : std_logic;
signal \un33_r_val_cry_7_THRU_CO\ : std_logic;
signal \N_95_cascade_\ : std_logic;
signal pwm_r_1_8 : std_logic;
signal \un34_r_val_0_cry_5_c_RNI0HHVZ0\ : std_logic;
signal \N_69_cascade_\ : std_logic;
signal \ctrZ0Z_26\ : std_logic;
signal pwm_b_1_6 : std_logic;
signal \ctrZ0Z_28\ : std_logic;
signal \pwm_r_1_cry_10_c_RNOZ0Z_0\ : std_logic;
signal pwm_r_1_10 : std_logic;
signal \un34_r_val_0_cry_3_c_RNIQ8FVZ0\ : std_logic;
signal \N_67_cascade_\ : std_logic;
signal pwm_b_1_4 : std_logic;
signal \ctrZ0Z_18\ : std_logic;
signal pwm_b_1_0 : std_logic;
signal \un34_r_val_0_cry_1_c_RNIK0DVZ0\ : std_logic;
signal \ctrZ0Z_20\ : std_logic;
signal \N_65_cascade_\ : std_logic;
signal pwm_b_1_2 : std_logic;
signal \ctrZ0Z_22\ : std_logic;
signal \ctrZ0Z_24\ : std_logic;
signal pwm_g_1_4 : std_logic;
signal pwm_g_1_7 : std_logic;
signal \un34_r_val_0_cry_6_c_RNI3LIVZ0\ : std_logic;
signal \ctrZ0Z_25\ : std_logic;
signal \ctrZ0Z_27\ : std_logic;
signal \ctrZ0Z_31\ : std_logic;
signal \N_70_cascade_\ : std_logic;
signal \ctrZ0Z_30\ : std_logic;
signal pwm_b_1_7 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \RGB1_wire\ : std_logic;
signal \RGB0_wire\ : std_logic;
signal \RGB2_wire\ : std_logic;

begin
    RGB1 <= \RGB1_wire\;
    RGB0 <= \RGB0_wire\;
    RGB2 <= \RGB2_wire\;

    \I__1133\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__4946\,
            I => pwm_b_1_4
        );

    \I__1131\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__4940\,
            I => \N__4935\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__4939\,
            I => \N__4932\
        );

    \I__1128\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4928\
        );

    \I__1127\ : Span4Mux_h
    port map (
            O => \N__4935\,
            I => \N__4925\
        );

    \I__1126\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4920\
        );

    \I__1125\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4920\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__4928\,
            I => \ctrZ0Z_18\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__4925\,
            I => \ctrZ0Z_18\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__4920\,
            I => \ctrZ0Z_18\
        );

    \I__1121\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4910\,
            I => pwm_b_1_0
        );

    \I__1119\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4903\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4900\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4896\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4893\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__4899\,
            I => \N__4890\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__4896\,
            I => \N__4885\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__4893\,
            I => \N__4885\
        );

    \I__1112\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4882\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__4885\,
            I => \un34_r_val_0_cry_1_c_RNIK0DVZ0\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__4882\,
            I => \un34_r_val_0_cry_1_c_RNIK0DVZ0\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__4877\,
            I => \N__4874\
        );

    \I__1108\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4869\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \N__4866\
        );

    \I__1106\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4862\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__4869\,
            I => \N__4859\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4856\
        );

    \I__1103\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4853\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4844\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__4859\,
            I => \N__4837\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__4856\,
            I => \N__4837\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__4853\,
            I => \N__4837\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4833\
        );

    \I__1097\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4822\
        );

    \I__1096\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4822\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4822\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4822\
        );

    \I__1093\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4822\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__4844\,
            I => \N__4817\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__4837\,
            I => \N__4817\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4814\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__4833\,
            I => \ctrZ0Z_20\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4822\,
            I => \ctrZ0Z_20\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__4817\,
            I => \ctrZ0Z_20\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__4814\,
            I => \ctrZ0Z_20\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__4805\,
            I => \N_65_cascade_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__4799\,
            I => pwm_b_1_2
        );

    \I__1082\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4790\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4785\
        );

    \I__1080\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4785\
        );

    \I__1079\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4781\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4790\,
            I => \N__4778\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__4785\,
            I => \N__4775\
        );

    \I__1076\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4772\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4781\,
            I => \N__4766\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__4778\,
            I => \N__4759\
        );

    \I__1073\ : Span4Mux_s2_v
    port map (
            O => \N__4775\,
            I => \N__4759\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4759\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \N__4755\
        );

    \I__1070\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4752\
        );

    \I__1069\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4749\
        );

    \I__1068\ : Span4Mux_h
    port map (
            O => \N__4766\,
            I => \N__4746\
        );

    \I__1067\ : Span4Mux_h
    port map (
            O => \N__4759\,
            I => \N__4743\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4738\
        );

    \I__1065\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4738\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4752\,
            I => \ctrZ0Z_22\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__4749\,
            I => \ctrZ0Z_22\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__4746\,
            I => \ctrZ0Z_22\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__4743\,
            I => \ctrZ0Z_22\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4738\,
            I => \ctrZ0Z_22\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4717\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4714\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4711\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4708\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4703\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4703\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \N__4699\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4696\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4693\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4684\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4684\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4708\,
            I => \N__4684\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4703\,
            I => \N__4684\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4679\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4679\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4696\,
            I => \N__4672\
        );

    \I__1043\ : Span4Mux_s2_v
    port map (
            O => \N__4693\,
            I => \N__4672\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__4684\,
            I => \N__4672\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__4679\,
            I => \N__4669\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__4672\,
            I => \ctrZ0Z_24\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__4669\,
            I => \ctrZ0Z_24\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__1035\ : Span4Mux_s3_h
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__4652\,
            I => pwm_g_1_4
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \N__4646\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__4637\,
            I => pwm_g_1_7
        );

    \I__1028\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4630\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4626\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4623\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__4629\,
            I => \N__4620\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4626\,
            I => \N__4617\
        );

    \I__1023\ : Span4Mux_h
    port map (
            O => \N__4623\,
            I => \N__4614\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4611\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__4617\,
            I => \un34_r_val_0_cry_6_c_RNI3LIVZ0\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__4614\,
            I => \un34_r_val_0_cry_6_c_RNI3LIVZ0\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4611\,
            I => \un34_r_val_0_cry_6_c_RNI3LIVZ0\
        );

    \I__1018\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4594\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4594\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4589\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4589\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__4600\,
            I => \N__4585\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4580\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4594\,
            I => \N__4577\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4589\,
            I => \N__4574\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4569\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4569\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4566\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4563\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4560\
        );

    \I__1005\ : Span4Mux_h
    port map (
            O => \N__4577\,
            I => \N__4557\
        );

    \I__1004\ : Span4Mux_h
    port map (
            O => \N__4574\,
            I => \N__4552\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4569\,
            I => \N__4552\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4566\,
            I => \ctrZ0Z_25\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4563\,
            I => \ctrZ0Z_25\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__4560\,
            I => \ctrZ0Z_25\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__4557\,
            I => \ctrZ0Z_25\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__4552\,
            I => \ctrZ0Z_25\
        );

    \I__997\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4536\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4529\
        );

    \I__995\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4525\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4522\
        );

    \I__993\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4517\
        );

    \I__992\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4517\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__4533\,
            I => \N__4514\
        );

    \I__990\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4509\
        );

    \I__989\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4509\
        );

    \I__988\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4505\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4498\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__4522\,
            I => \N__4498\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4498\
        );

    \I__984\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4495\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4509\,
            I => \N__4492\
        );

    \I__982\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4489\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4505\,
            I => \N__4484\
        );

    \I__980\ : Span4Mux_s2_v
    port map (
            O => \N__4498\,
            I => \N__4484\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4479\
        );

    \I__978\ : Span4Mux_v
    port map (
            O => \N__4492\,
            I => \N__4479\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4489\,
            I => \ctrZ0Z_27\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__4484\,
            I => \ctrZ0Z_27\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__4479\,
            I => \ctrZ0Z_27\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__973\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4453\
        );

    \I__972\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4453\
        );

    \I__971\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4448\
        );

    \I__970\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4448\
        );

    \I__969\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4443\
        );

    \I__968\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4443\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \N__4436\
        );

    \I__966\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4427\
        );

    \I__965\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4427\
        );

    \I__964\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4427\
        );

    \I__963\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4420\
        );

    \I__962\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4415\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4453\,
            I => \N__4407\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4448\,
            I => \N__4402\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4402\
        );

    \I__958\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4391\
        );

    \I__957\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4391\
        );

    \I__956\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4391\
        );

    \I__955\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4391\
        );

    \I__954\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4391\
        );

    \I__953\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4386\
        );

    \I__952\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4386\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4383\
        );

    \I__950\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4378\
        );

    \I__949\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4378\
        );

    \I__948\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4371\
        );

    \I__947\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4371\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4368\
        );

    \I__945\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4363\
        );

    \I__944\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4363\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4415\,
            I => \N__4358\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__4414\,
            I => \N__4354\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__4413\,
            I => \N__4350\
        );

    \I__940\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4341\
        );

    \I__939\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4341\
        );

    \I__938\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4341\
        );

    \I__937\ : Span4Mux_s3_v
    port map (
            O => \N__4407\,
            I => \N__4334\
        );

    \I__936\ : Span4Mux_s3_v
    port map (
            O => \N__4402\,
            I => \N__4334\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4391\,
            I => \N__4334\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4327\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__4383\,
            I => \N__4327\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4378\,
            I => \N__4327\
        );

    \I__931\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4324\
        );

    \I__930\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4321\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4371\,
            I => \N__4318\
        );

    \I__928\ : Span4Mux_s2_v
    port map (
            O => \N__4368\,
            I => \N__4313\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4363\,
            I => \N__4313\
        );

    \I__926\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4308\
        );

    \I__925\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4308\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__4358\,
            I => \N__4305\
        );

    \I__923\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4292\
        );

    \I__922\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4292\
        );

    \I__921\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4292\
        );

    \I__920\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4292\
        );

    \I__919\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4292\
        );

    \I__918\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4292\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4341\,
            I => \N__4287\
        );

    \I__916\ : Span4Mux_h
    port map (
            O => \N__4334\,
            I => \N__4287\
        );

    \I__915\ : Span4Mux_h
    port map (
            O => \N__4327\,
            I => \N__4284\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4324\,
            I => \ctrZ0Z_31\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4321\,
            I => \ctrZ0Z_31\
        );

    \I__912\ : Odrv4
    port map (
            O => \N__4318\,
            I => \ctrZ0Z_31\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__4313\,
            I => \ctrZ0Z_31\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4308\,
            I => \ctrZ0Z_31\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4305\,
            I => \ctrZ0Z_31\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4292\,
            I => \ctrZ0Z_31\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__4287\,
            I => \ctrZ0Z_31\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__4284\,
            I => \ctrZ0Z_31\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4265\,
            I => \N_70_cascade_\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4262\,
            I => \N__4250\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4261\,
            I => \N__4246\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__4260\,
            I => \N__4236\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__4259\,
            I => \N__4229\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \N__4218\
        );

    \I__899\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4210\
        );

    \I__898\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4210\
        );

    \I__897\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4210\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__4254\,
            I => \N__4206\
        );

    \I__895\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4190\
        );

    \I__894\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4190\
        );

    \I__893\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4190\
        );

    \I__892\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4190\
        );

    \I__891\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4190\
        );

    \I__890\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4190\
        );

    \I__889\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4190\
        );

    \I__888\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4177\
        );

    \I__887\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4177\
        );

    \I__886\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4177\
        );

    \I__885\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4177\
        );

    \I__884\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4177\
        );

    \I__883\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4177\
        );

    \I__882\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4164\
        );

    \I__881\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4164\
        );

    \I__880\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4164\
        );

    \I__879\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4164\
        );

    \I__878\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4164\
        );

    \I__877\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4164\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__4226\,
            I => \N__4156\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4225\,
            I => \N__4153\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__4224\,
            I => \N__4146\
        );

    \I__873\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4139\
        );

    \I__872\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4139\
        );

    \I__871\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4134\
        );

    \I__870\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4134\
        );

    \I__869\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4131\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4128\
        );

    \I__867\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4121\
        );

    \I__866\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4121\
        );

    \I__865\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4121\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4190\,
            I => \N__4114\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4177\,
            I => \N__4114\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4114\
        );

    \I__861\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4107\
        );

    \I__860\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4107\
        );

    \I__859\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4107\
        );

    \I__858\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4104\
        );

    \I__857\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4097\
        );

    \I__856\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4097\
        );

    \I__855\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4097\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__4152\,
            I => \N__4092\
        );

    \I__853\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4083\
        );

    \I__852\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4083\
        );

    \I__851\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4083\
        );

    \I__850\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4076\
        );

    \I__849\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4076\
        );

    \I__848\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4076\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4073\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4070\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4059\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__4128\,
            I => \N__4050\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4050\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__4114\,
            I => \N__4050\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4107\,
            I => \N__4050\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4104\,
            I => \N__4045\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4045\
        );

    \I__838\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4034\
        );

    \I__837\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4034\
        );

    \I__836\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4034\
        );

    \I__835\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4034\
        );

    \I__834\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4034\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4083\,
            I => \N__4025\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4076\,
            I => \N__4025\
        );

    \I__831\ : Span4Mux_h
    port map (
            O => \N__4073\,
            I => \N__4025\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__4070\,
            I => \N__4025\
        );

    \I__829\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4008\
        );

    \I__828\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4008\
        );

    \I__827\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4008\
        );

    \I__826\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4008\
        );

    \I__825\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4008\
        );

    \I__824\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4008\
        );

    \I__823\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4008\
        );

    \I__822\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4008\
        );

    \I__821\ : Span4Mux_h
    port map (
            O => \N__4059\,
            I => \N__4003\
        );

    \I__820\ : Span4Mux_h
    port map (
            O => \N__4050\,
            I => \N__4003\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__4045\,
            I => \ctrZ0Z_30\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4034\,
            I => \ctrZ0Z_30\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__4025\,
            I => \ctrZ0Z_30\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4008\,
            I => \ctrZ0Z_30\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__4003\,
            I => \ctrZ0Z_30\
        );

    \I__814\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3989\,
            I => pwm_b_1_7
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__3986\,
            I => \N__3982\
        );

    \I__811\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3978\
        );

    \I__810\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3975\
        );

    \I__809\ : InMux
    port map (
            O => \N__3981\,
            I => \N__3968\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3978\,
            I => \N__3965\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__3975\,
            I => \N__3962\
        );

    \I__806\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3957\
        );

    \I__805\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3957\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__3972\,
            I => \N__3953\
        );

    \I__803\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3949\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__3968\,
            I => \N__3946\
        );

    \I__801\ : Span4Mux_s2_v
    port map (
            O => \N__3965\,
            I => \N__3943\
        );

    \I__800\ : Span4Mux_h
    port map (
            O => \N__3962\,
            I => \N__3938\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__3957\,
            I => \N__3938\
        );

    \I__798\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3931\
        );

    \I__797\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3931\
        );

    \I__796\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3931\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3949\,
            I => \ctrZ0Z_29\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__3946\,
            I => \ctrZ0Z_29\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__3943\,
            I => \ctrZ0Z_29\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__3938\,
            I => \ctrZ0Z_29\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3931\,
            I => \ctrZ0Z_29\
        );

    \I__790\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3917\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3917\,
            I => \pwm_r_1_cry_11_c_RNOZ0Z_0\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__787\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3908\,
            I => pwm_r_1_11
        );

    \I__785\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__783\ : Span4Mux_s3_v
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__782\ : Odrv4
    port map (
            O => \N__3896\,
            I => pwm_g_1_6
        );

    \I__781\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__3890\,
            I => \N__3886\
        );

    \I__779\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3883\
        );

    \I__778\ : Span4Mux_s3_v
    port map (
            O => \N__3886\,
            I => \N__3877\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3883\,
            I => \N__3877\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__3882\,
            I => \N__3874\
        );

    \I__775\ : Span4Mux_h
    port map (
            O => \N__3877\,
            I => \N__3871\
        );

    \I__774\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3868\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__3871\,
            I => \un34_r_val_0_cry_7_c_RNI6PJVZ0\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__3868\,
            I => \un34_r_val_0_cry_7_c_RNI6PJVZ0\
        );

    \I__771\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3860\,
            I => \un33_r_val_cry_7_THRU_CO\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__3857\,
            I => \N_95_cascade_\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__767\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3848\,
            I => pwm_r_1_8
        );

    \I__765\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3842\,
            I => \N__3837\
        );

    \I__763\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3834\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__3840\,
            I => \N__3831\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__3837\,
            I => \N__3828\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3834\,
            I => \N__3825\
        );

    \I__759\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3822\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__3828\,
            I => \un34_r_val_0_cry_5_c_RNI0HHVZ0\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__3825\,
            I => \un34_r_val_0_cry_5_c_RNI0HHVZ0\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__3822\,
            I => \un34_r_val_0_cry_5_c_RNI0HHVZ0\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__3815\,
            I => \N_69_cascade_\
        );

    \I__754\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3808\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3811\,
            I => \N__3800\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3808\,
            I => \N__3797\
        );

    \I__751\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3790\
        );

    \I__750\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3790\
        );

    \I__749\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3790\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__3804\,
            I => \N__3786\
        );

    \I__747\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3782\
        );

    \I__746\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3779\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__3797\,
            I => \N__3774\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3790\,
            I => \N__3774\
        );

    \I__743\ : InMux
    port map (
            O => \N__3789\,
            I => \N__3769\
        );

    \I__742\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3769\
        );

    \I__741\ : InMux
    port map (
            O => \N__3785\,
            I => \N__3766\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3763\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3779\,
            I => \N__3758\
        );

    \I__738\ : Span4Mux_h
    port map (
            O => \N__3774\,
            I => \N__3758\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3769\,
            I => \N__3755\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3766\,
            I => \ctrZ0Z_26\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__3763\,
            I => \ctrZ0Z_26\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__3758\,
            I => \ctrZ0Z_26\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__3755\,
            I => \ctrZ0Z_26\
        );

    \I__732\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__3740\,
            I => pwm_b_1_6
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__3737\,
            I => \N__3732\
        );

    \I__728\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3725\
        );

    \I__727\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3725\
        );

    \I__726\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3719\
        );

    \I__725\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3713\
        );

    \I__724\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3713\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3725\,
            I => \N__3710\
        );

    \I__722\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3707\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__3723\,
            I => \N__3704\
        );

    \I__720\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3701\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3719\,
            I => \N__3698\
        );

    \I__718\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3695\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N__3692\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__3710\,
            I => \N__3687\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3707\,
            I => \N__3687\
        );

    \I__714\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3684\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3679\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__3698\,
            I => \N__3679\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3695\,
            I => \ctrZ0Z_28\
        );

    \I__710\ : Odrv4
    port map (
            O => \N__3692\,
            I => \ctrZ0Z_28\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__3687\,
            I => \ctrZ0Z_28\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3684\,
            I => \ctrZ0Z_28\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3679\,
            I => \ctrZ0Z_28\
        );

    \I__706\ : InMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3665\,
            I => \pwm_r_1_cry_10_c_RNOZ0Z_0\
        );

    \I__704\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3659\,
            I => pwm_r_1_10
        );

    \I__702\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3653\,
            I => \N__3649\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__3652\,
            I => \N__3645\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__3649\,
            I => \N__3642\
        );

    \I__698\ : InMux
    port map (
            O => \N__3648\,
            I => \N__3639\
        );

    \I__697\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3636\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__3642\,
            I => \un34_r_val_0_cry_3_c_RNIQ8FVZ0\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3639\,
            I => \un34_r_val_0_cry_3_c_RNIQ8FVZ0\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3636\,
            I => \un34_r_val_0_cry_3_c_RNIQ8FVZ0\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__3629\,
            I => \N_67_cascade_\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__691\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__3617\,
            I => pwm_r_1_2
        );

    \I__688\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3610\
        );

    \I__687\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3607\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3610\,
            I => \N__3600\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N__3600\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__3606\,
            I => \N__3592\
        );

    \I__683\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3589\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__3600\,
            I => \N__3586\
        );

    \I__681\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3583\
        );

    \I__680\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3576\
        );

    \I__679\ : InMux
    port map (
            O => \N__3597\,
            I => \N__3576\
        );

    \I__678\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3576\
        );

    \I__677\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3571\
        );

    \I__676\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3571\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3589\,
            I => \ctrZ0Z_21\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__3586\,
            I => \ctrZ0Z_21\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3583\,
            I => \ctrZ0Z_21\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3576\,
            I => \ctrZ0Z_21\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3571\,
            I => \ctrZ0Z_21\
        );

    \I__670\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3557\,
            I => \N__3552\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__3556\,
            I => \N__3549\
        );

    \I__667\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3546\
        );

    \I__666\ : Span4Mux_h
    port map (
            O => \N__3552\,
            I => \N__3543\
        );

    \I__665\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3540\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3546\,
            I => \un34_r_val_0_cry_2_c_RNIN4EVZ0\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__3543\,
            I => \un34_r_val_0_cry_2_c_RNIN4EVZ0\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3540\,
            I => \un34_r_val_0_cry_2_c_RNIN4EVZ0\
        );

    \I__661\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3530\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3530\,
            I => \un33_r_val_cry_2_THRU_CO\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__3527\,
            I => \N_90_cascade_\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__657\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3518\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3515\,
            I => pwm_r_1_3
        );

    \I__654\ : InMux
    port map (
            O => \N__3512\,
            I => \N__3509\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3509\,
            I => \un33_r_val_cry_5_THRU_CO\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__3506\,
            I => \N_93_cascade_\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__650\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3497\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3497\,
            I => pwm_r_1_6
        );

    \I__648\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3490\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__3493\,
            I => \N__3485\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3490\,
            I => \N__3482\
        );

    \I__645\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3479\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__3488\,
            I => \N__3474\
        );

    \I__643\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3469\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__3482\,
            I => \N__3464\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3464\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3478\,
            I => \N__3460\
        );

    \I__639\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3457\
        );

    \I__638\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3454\
        );

    \I__637\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3449\
        );

    \I__636\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3449\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3446\
        );

    \I__634\ : Span4Mux_h
    port map (
            O => \N__3464\,
            I => \N__3443\
        );

    \I__633\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3438\
        );

    \I__632\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3438\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3457\,
            I => \ctrZ0Z_23\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3454\,
            I => \ctrZ0Z_23\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3449\,
            I => \ctrZ0Z_23\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__3446\,
            I => \ctrZ0Z_23\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__3443\,
            I => \ctrZ0Z_23\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3438\,
            I => \ctrZ0Z_23\
        );

    \I__625\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3421\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__3424\,
            I => \N__3417\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3421\,
            I => \N__3414\
        );

    \I__622\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3411\
        );

    \I__621\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3408\
        );

    \I__620\ : Odrv4
    port map (
            O => \N__3414\,
            I => \un34_r_val_0_cry_4_c_RNITCGVZ0\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3411\,
            I => \un34_r_val_0_cry_4_c_RNITCGVZ0\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3408\,
            I => \un34_r_val_0_cry_4_c_RNITCGVZ0\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3401\,
            I => \N_68_cascade_\
        );

    \I__616\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3395\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3389\,
            I => pwm_b_1_5
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__611\ : InMux
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3380\,
            I => \un33_r_val_cry_6_THRU_CO\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \N_94_cascade_\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__607\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3368\,
            I => pwm_r_1_7
        );

    \I__605\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3362\,
            I => pwm_b_1_8
        );

    \I__603\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3355\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__3358\,
            I => \N__3352\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3348\
        );

    \I__600\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3345\
        );

    \I__599\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3342\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__3348\,
            I => pwm_ctr_i_8
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3345\,
            I => pwm_ctr_i_8
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3342\,
            I => pwm_ctr_i_8
        );

    \I__595\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3331\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \N__3328\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3331\,
            I => \N__3324\
        );

    \I__592\ : InMux
    port map (
            O => \N__3328\,
            I => \N__3321\
        );

    \I__591\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3318\
        );

    \I__590\ : Odrv4
    port map (
            O => \N__3324\,
            I => pwm_ctr_i_9
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3321\,
            I => pwm_ctr_i_9
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3318\,
            I => pwm_ctr_i_9
        );

    \I__587\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__585\ : Odrv12
    port map (
            O => \N__3305\,
            I => pwm_b_1_10
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__3302\,
            I => \N__3298\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__3301\,
            I => \N__3295\
        );

    \I__582\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3292\
        );

    \I__581\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3289\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3292\,
            I => \N__3285\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3289\,
            I => \N__3282\
        );

    \I__578\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3279\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__3285\,
            I => pwm_ctr_i_10
        );

    \I__576\ : Odrv4
    port map (
            O => \N__3282\,
            I => pwm_ctr_i_10
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3279\,
            I => pwm_ctr_i_10
        );

    \I__574\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__3266\,
            I => pwm_b_1_11
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__3263\,
            I => \N__3259\
        );

    \I__570\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3256\
        );

    \I__569\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3253\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3256\,
            I => \N__3249\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3253\,
            I => \N__3246\
        );

    \I__566\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3243\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__3249\,
            I => pwm_ctr_i_11
        );

    \I__564\ : Odrv4
    port map (
            O => \N__3246\,
            I => pwm_ctr_i_11
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3243\,
            I => pwm_ctr_i_11
        );

    \I__562\ : InMux
    port map (
            O => \N__3236\,
            I => pwm_b_1
        );

    \I__561\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__3227\,
            I => \pwm_bZ0\
        );

    \I__558\ : ClkMux
    port map (
            O => \N__3224\,
            I => \N__3197\
        );

    \I__557\ : ClkMux
    port map (
            O => \N__3223\,
            I => \N__3197\
        );

    \I__556\ : ClkMux
    port map (
            O => \N__3222\,
            I => \N__3197\
        );

    \I__555\ : ClkMux
    port map (
            O => \N__3221\,
            I => \N__3197\
        );

    \I__554\ : ClkMux
    port map (
            O => \N__3220\,
            I => \N__3197\
        );

    \I__553\ : ClkMux
    port map (
            O => \N__3219\,
            I => \N__3197\
        );

    \I__552\ : ClkMux
    port map (
            O => \N__3218\,
            I => \N__3197\
        );

    \I__551\ : ClkMux
    port map (
            O => \N__3217\,
            I => \N__3197\
        );

    \I__550\ : ClkMux
    port map (
            O => \N__3216\,
            I => \N__3197\
        );

    \I__549\ : GlobalMux
    port map (
            O => \N__3197\,
            I => clk
        );

    \I__548\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3191\,
            I => \N__3187\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__3190\,
            I => \N__3183\
        );

    \I__545\ : Span4Mux_s1_v
    port map (
            O => \N__3187\,
            I => \N__3180\
        );

    \I__544\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3177\
        );

    \I__543\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3174\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__3180\,
            I => \un34_r_val_0_cry_8_c_RNI9TKVZ0\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3177\,
            I => \un34_r_val_0_cry_8_c_RNI9TKVZ0\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3174\,
            I => \un34_r_val_0_cry_8_c_RNI9TKVZ0\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__3167\,
            I => \N_72_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3161\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3161\,
            I => pwm_b_1_9
        );

    \I__536\ : InMux
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3155\,
            I => \un33_r_val_cry_1_THRU_CO\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3152\,
            I => \N_89_cascade_\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3149\,
            I => \N__3145\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__531\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3138\
        );

    \I__530\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3135\
        );

    \I__529\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3132\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3138\,
            I => \N__3129\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3135\,
            I => pwm_ctr_i_0
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3132\,
            I => pwm_ctr_i_0
        );

    \I__525\ : Odrv4
    port map (
            O => \N__3129\,
            I => pwm_ctr_i_0
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3122\,
            I => \N__3118\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3121\,
            I => \N__3115\
        );

    \I__522\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3112\
        );

    \I__521\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3108\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3112\,
            I => \N__3105\
        );

    \I__519\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3102\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3108\,
            I => \N__3097\
        );

    \I__517\ : Span4Mux_h
    port map (
            O => \N__3105\,
            I => \N__3097\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3102\,
            I => pwm_ctr_i_1
        );

    \I__515\ : Odrv4
    port map (
            O => \N__3097\,
            I => pwm_ctr_i_1
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__513\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3086\,
            I => pwm_b_1_1
        );

    \I__511\ : InMux
    port map (
            O => \N__3083\,
            I => \N__3079\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \N__3076\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3079\,
            I => \N__3072\
        );

    \I__508\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3069\
        );

    \I__507\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3066\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3072\,
            I => pwm_ctr_i_2
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3069\,
            I => pwm_ctr_i_2
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3066\,
            I => pwm_ctr_i_2
        );

    \I__503\ : InMux
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__3053\,
            I => pwm_b_1_3
        );

    \I__500\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3046\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__3049\,
            I => \N__3043\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3046\,
            I => \N__3039\
        );

    \I__497\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3036\
        );

    \I__496\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3033\
        );

    \I__495\ : Odrv4
    port map (
            O => \N__3039\,
            I => pwm_ctr_i_3
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3036\,
            I => pwm_ctr_i_3
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3033\,
            I => pwm_ctr_i_3
        );

    \I__492\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3023\,
            I => \N__3019\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3022\,
            I => \N__3016\
        );

    \I__489\ : Span4Mux_h
    port map (
            O => \N__3019\,
            I => \N__3012\
        );

    \I__488\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3009\
        );

    \I__487\ : InMux
    port map (
            O => \N__3015\,
            I => \N__3006\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__3012\,
            I => pwm_ctr_i_4
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3009\,
            I => pwm_ctr_i_4
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3006\,
            I => pwm_ctr_i_4
        );

    \I__483\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2995\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__2998\,
            I => \N__2992\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2995\,
            I => \N__2988\
        );

    \I__480\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2985\
        );

    \I__479\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2982\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__2988\,
            I => pwm_ctr_i_5
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2985\,
            I => pwm_ctr_i_5
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2982\,
            I => pwm_ctr_i_5
        );

    \I__475\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2970\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__2974\,
            I => \N__2967\
        );

    \I__473\ : CascadeMux
    port map (
            O => \N__2973\,
            I => \N__2964\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2970\,
            I => \N__2961\
        );

    \I__471\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2958\
        );

    \I__470\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2955\
        );

    \I__469\ : Span4Mux_h
    port map (
            O => \N__2961\,
            I => \N__2952\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2958\,
            I => pwm_ctr_i_6
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2955\,
            I => pwm_ctr_i_6
        );

    \I__466\ : Odrv4
    port map (
            O => \N__2952\,
            I => pwm_ctr_i_6
        );

    \I__465\ : InMux
    port map (
            O => \N__2945\,
            I => \N__2941\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2941\,
            I => \N__2935\
        );

    \I__462\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2932\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__2935\,
            I => \N__2928\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2932\,
            I => \N__2925\
        );

    \I__459\ : InMux
    port map (
            O => \N__2931\,
            I => \N__2922\
        );

    \I__458\ : Odrv4
    port map (
            O => \N__2928\,
            I => pwm_ctr_i_7
        );

    \I__457\ : Odrv4
    port map (
            O => \N__2925\,
            I => pwm_ctr_i_7
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2922\,
            I => pwm_ctr_i_7
        );

    \I__455\ : InMux
    port map (
            O => \N__2915\,
            I => pwm_r_1
        );

    \I__454\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__452\ : Span4Mux_s2_v
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__451\ : Odrv4
    port map (
            O => \N__2903\,
            I => \pwm_rZ0\
        );

    \I__450\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2894\,
            I => \un33_r_val_cry_8_THRU_CO\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__2891\,
            I => \N_96_cascade_\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__445\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2882\,
            I => pwm_r_1_9
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__2879\,
            I => \N__2875\
        );

    \I__442\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__441\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2872\,
            I => \un34_r_val_0_cry_9_c_RNIV0HKZ0\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2869\,
            I => \un34_r_val_0_cry_9_c_RNIV0HKZ0\
        );

    \I__438\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2861\,
            I => \un33_r_val_cry_3_THRU_CO\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__2858\,
            I => \N_91_cascade_\
        );

    \I__435\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2852\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2852\,
            I => pwm_r_1_0
        );

    \I__433\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__2843\,
            I => pwm_r_1_1
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__2840\,
            I => \N__2837\
        );

    \I__429\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2834\,
            I => pwm_r_1_4
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__426\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2825\,
            I => pwm_r_1_5
        );

    \I__424\ : InMux
    port map (
            O => \N__2822\,
            I => un33_r_val_cry_3
        );

    \I__423\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__2813\,
            I => \un33_r_val_cry_4_THRU_CO\
        );

    \I__420\ : InMux
    port map (
            O => \N__2810\,
            I => un33_r_val_cry_4
        );

    \I__419\ : InMux
    port map (
            O => \N__2807\,
            I => un33_r_val_cry_5
        );

    \I__418\ : InMux
    port map (
            O => \N__2804\,
            I => un33_r_val_cry_6
        );

    \I__417\ : InMux
    port map (
            O => \N__2801\,
            I => \bfn_3_26_0_\
        );

    \I__416\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2791\
        );

    \I__414\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2787\
        );

    \I__413\ : Span4Mux_v
    port map (
            O => \N__2791\,
            I => \N__2783\
        );

    \I__412\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2780\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2787\,
            I => \N__2777\
        );

    \I__410\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2774\
        );

    \I__409\ : Sp12to4
    port map (
            O => \N__2783\,
            I => \N__2770\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2780\,
            I => \N__2763\
        );

    \I__407\ : Span4Mux_s1_v
    port map (
            O => \N__2777\,
            I => \N__2763\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2774\,
            I => \N__2763\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__2773\,
            I => \N__2752\
        );

    \I__404\ : Span12Mux_h
    port map (
            O => \N__2770\,
            I => \N__2749\
        );

    \I__403\ : Span4Mux_v
    port map (
            O => \N__2763\,
            I => \N__2746\
        );

    \I__402\ : InMux
    port map (
            O => \N__2762\,
            I => \N__2743\
        );

    \I__401\ : InMux
    port map (
            O => \N__2761\,
            I => \N__2740\
        );

    \I__400\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2733\
        );

    \I__399\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2733\
        );

    \I__398\ : InMux
    port map (
            O => \N__2758\,
            I => \N__2733\
        );

    \I__397\ : InMux
    port map (
            O => \N__2757\,
            I => \N__2724\
        );

    \I__396\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2724\
        );

    \I__395\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2724\
        );

    \I__394\ : InMux
    port map (
            O => \N__2752\,
            I => \N__2724\
        );

    \I__393\ : Odrv12
    port map (
            O => \N__2749\,
            I => \CONSTANT_ONE_NET\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__2746\,
            I => \CONSTANT_ONE_NET\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2743\,
            I => \CONSTANT_ONE_NET\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2740\,
            I => \CONSTANT_ONE_NET\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2733\,
            I => \CONSTANT_ONE_NET\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2724\,
            I => \CONSTANT_ONE_NET\
        );

    \I__387\ : InMux
    port map (
            O => \N__2711\,
            I => un33_r_val_cry_8
        );

    \I__386\ : InMux
    port map (
            O => \N__2708\,
            I => un33_r_val_cry_9
        );

    \I__385\ : InMux
    port map (
            O => \N__2705\,
            I => un33_r_val_cry_10
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__2702\,
            I => \un33_r_val_cry_10_THRU_CO_cascade_\
        );

    \I__383\ : InMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2696\,
            I => \un34_r_val_0_cry_10_THRU_CO\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__380\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__2684\,
            I => pwm_g_1_11
        );

    \I__377\ : InMux
    port map (
            O => \N__2681\,
            I => pwm_g_1
        );

    \I__376\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2675\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2675\,
            I => \N__2672\
        );

    \I__374\ : Odrv4
    port map (
            O => \N__2672\,
            I => \pwm_gZ0\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__2669\,
            I => \N_71_cascade_\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__2666\,
            I => \N__2663\
        );

    \I__371\ : InMux
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2660\,
            I => pwm_g_1_10
        );

    \I__369\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2653\
        );

    \I__368\ : InMux
    port map (
            O => \N__2656\,
            I => \N__2650\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2653\,
            I => \ctr_RNI7D9MZ0Z_21\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2650\,
            I => \ctr_RNI7D9MZ0Z_21\
        );

    \I__365\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2642\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2642\,
            I => \un33_r_val_cry_0_THRU_CO\
        );

    \I__363\ : InMux
    port map (
            O => \N__2639\,
            I => un33_r_val_cry_0
        );

    \I__362\ : InMux
    port map (
            O => \N__2636\,
            I => un33_r_val_cry_1
        );

    \I__361\ : InMux
    port map (
            O => \N__2633\,
            I => un33_r_val_cry_2
        );

    \I__360\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2626\
        );

    \I__359\ : InMux
    port map (
            O => \N__2629\,
            I => \N__2623\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2626\,
            I => \pwm_ctrZ0Z_3\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2623\,
            I => \pwm_ctrZ0Z_3\
        );

    \I__356\ : CascadeMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__355\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2612\,
            I => pwm_g_1_3
        );

    \I__353\ : InMux
    port map (
            O => \N__2609\,
            I => \N__2605\
        );

    \I__352\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2602\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2605\,
            I => \pwm_ctrZ0Z_4\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2602\,
            I => \pwm_ctrZ0Z_4\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__348\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__346\ : Span4Mux_s2_v
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__2585\,
            I => pwm_g_1_5
        );

    \I__344\ : InMux
    port map (
            O => \N__2582\,
            I => \N__2578\
        );

    \I__343\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2575\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2578\,
            I => \pwm_ctrZ0Z_5\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2575\,
            I => \pwm_ctrZ0Z_5\
        );

    \I__340\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2566\
        );

    \I__339\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2563\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2566\,
            I => \pwm_ctrZ0Z_6\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2563\,
            I => \pwm_ctrZ0Z_6\
        );

    \I__336\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2554\
        );

    \I__335\ : InMux
    port map (
            O => \N__2557\,
            I => \N__2551\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2554\,
            I => \pwm_ctrZ0Z_7\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2551\,
            I => \pwm_ctrZ0Z_7\
        );

    \I__332\ : CascadeMux
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__331\ : InMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2540\,
            I => pwm_g_1_8
        );

    \I__329\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2533\
        );

    \I__328\ : InMux
    port map (
            O => \N__2536\,
            I => \N__2530\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2533\,
            I => \pwm_ctrZ0Z_8\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2530\,
            I => \pwm_ctrZ0Z_8\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__324\ : InMux
    port map (
            O => \N__2522\,
            I => \N__2519\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__322\ : Odrv4
    port map (
            O => \N__2516\,
            I => pwm_g_1_9
        );

    \I__321\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2509\
        );

    \I__320\ : InMux
    port map (
            O => \N__2512\,
            I => \N__2506\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2509\,
            I => \pwm_ctrZ0Z_9\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2506\,
            I => \pwm_ctrZ0Z_9\
        );

    \I__317\ : InMux
    port map (
            O => \N__2501\,
            I => \N__2497\
        );

    \I__316\ : InMux
    port map (
            O => \N__2500\,
            I => \N__2494\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2497\,
            I => \pwm_ctrZ0Z_10\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2494\,
            I => \pwm_ctrZ0Z_10\
        );

    \I__313\ : InMux
    port map (
            O => \N__2489\,
            I => \N__2485\
        );

    \I__312\ : InMux
    port map (
            O => \N__2488\,
            I => \N__2482\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2485\,
            I => \pwm_ctrZ0Z_11\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2482\,
            I => \pwm_ctrZ0Z_11\
        );

    \I__309\ : CascadeMux
    port map (
            O => \N__2477\,
            I => \N_87_cascade_\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2474\,
            I => \N__2471\
        );

    \I__307\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2468\,
            I => \N__2462\
        );

    \I__305\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2459\
        );

    \I__304\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2454\
        );

    \I__303\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2454\
        );

    \I__302\ : Span4Mux_v
    port map (
            O => \N__2462\,
            I => \N__2451\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2459\,
            I => \ctrZ0Z_19\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2454\,
            I => \ctrZ0Z_19\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__2451\,
            I => \ctrZ0Z_19\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__2444\,
            I => \un40_b_val_3_ns_1_1_cascade_\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2441\,
            I => \N__2438\
        );

    \I__296\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2435\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2435\,
            I => pwm_g_1_0
        );

    \I__294\ : InMux
    port map (
            O => \N__2432\,
            I => \N__2428\
        );

    \I__293\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2425\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2428\,
            I => \pwm_ctrZ0Z_0\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2425\,
            I => \pwm_ctrZ0Z_0\
        );

    \I__290\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2416\
        );

    \I__289\ : InMux
    port map (
            O => \N__2419\,
            I => \N__2413\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2416\,
            I => \pwm_ctrZ0Z_1\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2413\,
            I => \pwm_ctrZ0Z_1\
        );

    \I__286\ : InMux
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2405\,
            I => pwm_g_1_1
        );

    \I__284\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2398\
        );

    \I__283\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2395\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2398\,
            I => \pwm_ctrZ0Z_2\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2395\,
            I => \pwm_ctrZ0Z_2\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__279\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2384\,
            I => pwm_g_1_2
        );

    \I__277\ : InMux
    port map (
            O => \N__2381\,
            I => un34_r_val_0_cry_9
        );

    \I__276\ : InMux
    port map (
            O => \N__2378\,
            I => un34_r_val_0_cry_10
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__2375\,
            I => \un34_r_val_0_cry_10_THRU_CO_cascade_\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2372\,
            I => \N_92_cascade_\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2369\,
            I => \N_66_cascade_\
        );

    \I__272\ : InMux
    port map (
            O => \N__2366\,
            I => un34_r_val_0_cry_1
        );

    \I__271\ : InMux
    port map (
            O => \N__2363\,
            I => un34_r_val_0_cry_2
        );

    \I__270\ : InMux
    port map (
            O => \N__2360\,
            I => un34_r_val_0_cry_3
        );

    \I__269\ : InMux
    port map (
            O => \N__2357\,
            I => un34_r_val_0_cry_4
        );

    \I__268\ : InMux
    port map (
            O => \N__2354\,
            I => un34_r_val_0_cry_5
        );

    \I__267\ : InMux
    port map (
            O => \N__2351\,
            I => un34_r_val_0_cry_6
        );

    \I__266\ : InMux
    port map (
            O => \N__2348\,
            I => un34_r_val_0_cry_7
        );

    \I__265\ : InMux
    port map (
            O => \N__2345\,
            I => \bfn_2_27_0_\
        );

    \I__264\ : InMux
    port map (
            O => \N__2342\,
            I => pwm_ctr_cry_8
        );

    \I__263\ : InMux
    port map (
            O => \N__2339\,
            I => pwm_ctr_cry_9
        );

    \I__262\ : InMux
    port map (
            O => \N__2336\,
            I => pwm_ctr_cry_10
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__2333\,
            I => \N_88_cascade_\
        );

    \I__260\ : InMux
    port map (
            O => \N__2330\,
            I => \bfn_1_29_0_\
        );

    \I__259\ : InMux
    port map (
            O => \N__2327\,
            I => pwm_ctr_cry_0
        );

    \I__258\ : InMux
    port map (
            O => \N__2324\,
            I => pwm_ctr_cry_1
        );

    \I__257\ : InMux
    port map (
            O => \N__2321\,
            I => pwm_ctr_cry_2
        );

    \I__256\ : InMux
    port map (
            O => \N__2318\,
            I => pwm_ctr_cry_3
        );

    \I__255\ : InMux
    port map (
            O => \N__2315\,
            I => pwm_ctr_cry_4
        );

    \I__254\ : InMux
    port map (
            O => \N__2312\,
            I => pwm_ctr_cry_5
        );

    \I__253\ : InMux
    port map (
            O => \N__2309\,
            I => pwm_ctr_cry_6
        );

    \I__252\ : InMux
    port map (
            O => \N__2306\,
            I => \bfn_1_30_0_\
        );

    \I__251\ : InMux
    port map (
            O => \N__2303\,
            I => ctr_cry_22
        );

    \I__250\ : InMux
    port map (
            O => \N__2300\,
            I => \bfn_1_28_0_\
        );

    \I__249\ : InMux
    port map (
            O => \N__2297\,
            I => ctr_cry_24
        );

    \I__248\ : InMux
    port map (
            O => \N__2294\,
            I => ctr_cry_25
        );

    \I__247\ : InMux
    port map (
            O => \N__2291\,
            I => ctr_cry_26
        );

    \I__246\ : InMux
    port map (
            O => \N__2288\,
            I => ctr_cry_27
        );

    \I__245\ : InMux
    port map (
            O => \N__2285\,
            I => ctr_cry_28
        );

    \I__244\ : InMux
    port map (
            O => \N__2282\,
            I => ctr_cry_29
        );

    \I__243\ : InMux
    port map (
            O => \N__2279\,
            I => ctr_cry_30
        );

    \I__242\ : InMux
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2273\,
            I => \ctrZ0Z_14\
        );

    \I__240\ : InMux
    port map (
            O => \N__2270\,
            I => ctr_cry_13
        );

    \I__239\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2264\,
            I => \ctrZ0Z_15\
        );

    \I__237\ : InMux
    port map (
            O => \N__2261\,
            I => ctr_cry_14
        );

    \I__236\ : InMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2255\,
            I => \ctrZ0Z_16\
        );

    \I__234\ : InMux
    port map (
            O => \N__2252\,
            I => \bfn_1_27_0_\
        );

    \I__233\ : InMux
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2246\,
            I => \ctrZ0Z_17\
        );

    \I__231\ : InMux
    port map (
            O => \N__2243\,
            I => ctr_cry_16
        );

    \I__230\ : InMux
    port map (
            O => \N__2240\,
            I => ctr_cry_17
        );

    \I__229\ : InMux
    port map (
            O => \N__2237\,
            I => ctr_cry_18
        );

    \I__228\ : InMux
    port map (
            O => \N__2234\,
            I => ctr_cry_19
        );

    \I__227\ : InMux
    port map (
            O => \N__2231\,
            I => ctr_cry_20
        );

    \I__226\ : InMux
    port map (
            O => \N__2228\,
            I => ctr_cry_21
        );

    \I__225\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2222\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2222\,
            I => \ctrZ0Z_6\
        );

    \I__223\ : InMux
    port map (
            O => \N__2219\,
            I => ctr_cry_5
        );

    \I__222\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2213\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2213\,
            I => \ctrZ0Z_7\
        );

    \I__220\ : InMux
    port map (
            O => \N__2210\,
            I => ctr_cry_6
        );

    \I__219\ : InMux
    port map (
            O => \N__2207\,
            I => \N__2204\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2204\,
            I => \ctrZ0Z_8\
        );

    \I__217\ : InMux
    port map (
            O => \N__2201\,
            I => \bfn_1_26_0_\
        );

    \I__216\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2195\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2195\,
            I => \ctrZ0Z_9\
        );

    \I__214\ : InMux
    port map (
            O => \N__2192\,
            I => ctr_cry_8
        );

    \I__213\ : InMux
    port map (
            O => \N__2189\,
            I => \N__2186\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2186\,
            I => \ctrZ0Z_10\
        );

    \I__211\ : InMux
    port map (
            O => \N__2183\,
            I => ctr_cry_9
        );

    \I__210\ : InMux
    port map (
            O => \N__2180\,
            I => \N__2177\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__2177\,
            I => \ctrZ0Z_11\
        );

    \I__208\ : InMux
    port map (
            O => \N__2174\,
            I => ctr_cry_10
        );

    \I__207\ : InMux
    port map (
            O => \N__2171\,
            I => \N__2168\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__2168\,
            I => \ctrZ0Z_12\
        );

    \I__205\ : InMux
    port map (
            O => \N__2165\,
            I => ctr_cry_11
        );

    \I__204\ : InMux
    port map (
            O => \N__2162\,
            I => \N__2159\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__2159\,
            I => \ctrZ0Z_13\
        );

    \I__202\ : InMux
    port map (
            O => \N__2156\,
            I => ctr_cry_12
        );

    \I__201\ : InMux
    port map (
            O => \N__2153\,
            I => \N__2150\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2150\,
            I => \ctrZ0Z_0\
        );

    \I__199\ : InMux
    port map (
            O => \N__2147\,
            I => \bfn_1_25_0_\
        );

    \I__198\ : InMux
    port map (
            O => \N__2144\,
            I => \N__2141\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2141\,
            I => \ctrZ0Z_1\
        );

    \I__196\ : InMux
    port map (
            O => \N__2138\,
            I => ctr_cry_0
        );

    \I__195\ : InMux
    port map (
            O => \N__2135\,
            I => \N__2132\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__2132\,
            I => \ctrZ0Z_2\
        );

    \I__193\ : InMux
    port map (
            O => \N__2129\,
            I => ctr_cry_1
        );

    \I__192\ : InMux
    port map (
            O => \N__2126\,
            I => \N__2123\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__2123\,
            I => \ctrZ0Z_3\
        );

    \I__190\ : InMux
    port map (
            O => \N__2120\,
            I => ctr_cry_2
        );

    \I__189\ : InMux
    port map (
            O => \N__2117\,
            I => \N__2114\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__2114\,
            I => \ctrZ0Z_4\
        );

    \I__187\ : InMux
    port map (
            O => \N__2111\,
            I => ctr_cry_3
        );

    \I__186\ : InMux
    port map (
            O => \N__2108\,
            I => \N__2105\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__2105\,
            I => \ctrZ0Z_5\
        );

    \I__184\ : InMux
    port map (
            O => \N__2102\,
            I => ctr_cry_4
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un33_r_val_cry_7,
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_3_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_27_0_\
        );

    \IN_MUX_bfv_3_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => pwm_r_1_cry_7,
            carryinitout => \bfn_3_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_3_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => pwm_b_1_cry_7,
            carryinitout => \bfn_3_30_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => pwm_g_1_cry_7,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => pwm_ctr_cry_7,
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => ctr_cry_7,
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_1_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => ctr_cry_15,
            carryinitout => \bfn_1_27_0_\
        );

    \IN_MUX_bfv_1_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => ctr_cry_23,
            carryinitout => \bfn_1_28_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un34_r_val_0_cry_8,
            carryinitout => \bfn_2_27_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \RGBA_DRIVER\ : SB_RGBA_DRV
    generic map (
            CURRENT_MODE => "0b1",
            RGB2_CURRENT => "0b000111",
            RGB1_CURRENT => "0b000111",
            RGB0_CURRENT => "0b000111"
        )
    port map (
            RGBLEDEN => \N__2794\,
            RGB2PWM => \N__2912\,
            RGB1 => \RGB1_wire\,
            CURREN => \N__2798\,
            RGB2 => \RGB2_wire\,
            RGB1PWM => \N__3233\,
            RGB0PWM => \N__2678\,
            RGB0 => \RGB0_wire\
        );

    \inthosc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b00"
        )
    port map (
            CLKHFPU => \N__2786\,
            CLKHFEN => \N__2790\,
            CLKHF => clk
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \ctr_0_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2153\,
            in2 => \_gnd_net_\,
            in3 => \N__2147\,
            lcout => \ctrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => ctr_cry_0,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_1_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2144\,
            in2 => \_gnd_net_\,
            in3 => \N__2138\,
            lcout => \ctrZ0Z_1\,
            ltout => OPEN,
            carryin => ctr_cry_0,
            carryout => ctr_cry_1,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_2_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2135\,
            in2 => \_gnd_net_\,
            in3 => \N__2129\,
            lcout => \ctrZ0Z_2\,
            ltout => OPEN,
            carryin => ctr_cry_1,
            carryout => ctr_cry_2,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_3_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2126\,
            in2 => \_gnd_net_\,
            in3 => \N__2120\,
            lcout => \ctrZ0Z_3\,
            ltout => OPEN,
            carryin => ctr_cry_2,
            carryout => ctr_cry_3,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_4_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2117\,
            in2 => \_gnd_net_\,
            in3 => \N__2111\,
            lcout => \ctrZ0Z_4\,
            ltout => OPEN,
            carryin => ctr_cry_3,
            carryout => ctr_cry_4,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_5_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2108\,
            in2 => \_gnd_net_\,
            in3 => \N__2102\,
            lcout => \ctrZ0Z_5\,
            ltout => OPEN,
            carryin => ctr_cry_4,
            carryout => ctr_cry_5,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_6_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2225\,
            in2 => \_gnd_net_\,
            in3 => \N__2219\,
            lcout => \ctrZ0Z_6\,
            ltout => OPEN,
            carryin => ctr_cry_5,
            carryout => ctr_cry_6,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_7_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2216\,
            in2 => \_gnd_net_\,
            in3 => \N__2210\,
            lcout => \ctrZ0Z_7\,
            ltout => OPEN,
            carryin => ctr_cry_6,
            carryout => ctr_cry_7,
            clk => \N__3224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_8_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2207\,
            in2 => \_gnd_net_\,
            in3 => \N__2201\,
            lcout => \ctrZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => ctr_cry_8,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_9_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2198\,
            in2 => \_gnd_net_\,
            in3 => \N__2192\,
            lcout => \ctrZ0Z_9\,
            ltout => OPEN,
            carryin => ctr_cry_8,
            carryout => ctr_cry_9,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_10_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2189\,
            in2 => \_gnd_net_\,
            in3 => \N__2183\,
            lcout => \ctrZ0Z_10\,
            ltout => OPEN,
            carryin => ctr_cry_9,
            carryout => ctr_cry_10,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_11_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2180\,
            in2 => \_gnd_net_\,
            in3 => \N__2174\,
            lcout => \ctrZ0Z_11\,
            ltout => OPEN,
            carryin => ctr_cry_10,
            carryout => ctr_cry_11,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_12_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2171\,
            in2 => \_gnd_net_\,
            in3 => \N__2165\,
            lcout => \ctrZ0Z_12\,
            ltout => OPEN,
            carryin => ctr_cry_11,
            carryout => ctr_cry_12,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_13_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2162\,
            in2 => \_gnd_net_\,
            in3 => \N__2156\,
            lcout => \ctrZ0Z_13\,
            ltout => OPEN,
            carryin => ctr_cry_12,
            carryout => ctr_cry_13,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_14_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2276\,
            in2 => \_gnd_net_\,
            in3 => \N__2270\,
            lcout => \ctrZ0Z_14\,
            ltout => OPEN,
            carryin => ctr_cry_13,
            carryout => ctr_cry_14,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_15_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2267\,
            in2 => \_gnd_net_\,
            in3 => \N__2261\,
            lcout => \ctrZ0Z_15\,
            ltout => OPEN,
            carryin => ctr_cry_14,
            carryout => ctr_cry_15,
            clk => \N__3222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_16_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2258\,
            in2 => \_gnd_net_\,
            in3 => \N__2252\,
            lcout => \ctrZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_27_0_\,
            carryout => ctr_cry_16,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_17_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2249\,
            in2 => \_gnd_net_\,
            in3 => \N__2243\,
            lcout => \ctrZ0Z_17\,
            ltout => OPEN,
            carryin => ctr_cry_16,
            carryout => ctr_cry_17,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_18_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4938\,
            in2 => \_gnd_net_\,
            in3 => \N__2240\,
            lcout => \ctrZ0Z_18\,
            ltout => OPEN,
            carryin => ctr_cry_17,
            carryout => ctr_cry_18,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_19_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2467\,
            in2 => \_gnd_net_\,
            in3 => \N__2237\,
            lcout => \ctrZ0Z_19\,
            ltout => OPEN,
            carryin => ctr_cry_18,
            carryout => ctr_cry_19,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_20_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4852\,
            in2 => \_gnd_net_\,
            in3 => \N__2234\,
            lcout => \ctrZ0Z_20\,
            ltout => OPEN,
            carryin => ctr_cry_19,
            carryout => ctr_cry_20,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_21_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__2231\,
            lcout => \ctrZ0Z_21\,
            ltout => OPEN,
            carryin => ctr_cry_20,
            carryout => ctr_cry_21,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_22_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4770\,
            in2 => \_gnd_net_\,
            in3 => \N__2228\,
            lcout => \ctrZ0Z_22\,
            ltout => OPEN,
            carryin => ctr_cry_21,
            carryout => ctr_cry_22,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_23_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3477\,
            in2 => \_gnd_net_\,
            in3 => \N__2303\,
            lcout => \ctrZ0Z_23\,
            ltout => OPEN,
            carryin => ctr_cry_22,
            carryout => ctr_cry_23,
            clk => \N__3221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_24_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4720\,
            in2 => \_gnd_net_\,
            in3 => \N__2300\,
            lcout => \ctrZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_1_28_0_\,
            carryout => ctr_cry_24,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_25_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4584\,
            in2 => \_gnd_net_\,
            in3 => \N__2297\,
            lcout => \ctrZ0Z_25\,
            ltout => OPEN,
            carryin => ctr_cry_24,
            carryout => ctr_cry_25,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_26_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3785\,
            in2 => \_gnd_net_\,
            in3 => \N__2294\,
            lcout => \ctrZ0Z_26\,
            ltout => OPEN,
            carryin => ctr_cry_25,
            carryout => ctr_cry_26,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_27_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4508\,
            in2 => \_gnd_net_\,
            in3 => \N__2291\,
            lcout => \ctrZ0Z_27\,
            ltout => OPEN,
            carryin => ctr_cry_26,
            carryout => ctr_cry_27,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_28_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3718\,
            in2 => \_gnd_net_\,
            in3 => \N__2288\,
            lcout => \ctrZ0Z_28\,
            ltout => OPEN,
            carryin => ctr_cry_27,
            carryout => ctr_cry_28,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_29_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3971\,
            in2 => \_gnd_net_\,
            in3 => \N__2285\,
            lcout => \ctrZ0Z_29\,
            ltout => OPEN,
            carryin => ctr_cry_28,
            carryout => ctr_cry_29,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_30_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4160\,
            in2 => \_gnd_net_\,
            in3 => \N__2282\,
            lcout => \ctrZ0Z_30\,
            ltout => OPEN,
            carryin => ctr_cry_29,
            carryout => ctr_cry_30,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_31_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4377\,
            in2 => \_gnd_net_\,
            in3 => \N__2279\,
            lcout => \ctrZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_0_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2432\,
            in2 => \_gnd_net_\,
            in3 => \N__2330\,
            lcout => \pwm_ctrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => pwm_ctr_cry_0,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_1_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2420\,
            in2 => \_gnd_net_\,
            in3 => \N__2327\,
            lcout => \pwm_ctrZ0Z_1\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_0,
            carryout => pwm_ctr_cry_1,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_2_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2402\,
            in2 => \_gnd_net_\,
            in3 => \N__2324\,
            lcout => \pwm_ctrZ0Z_2\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_1,
            carryout => pwm_ctr_cry_2,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_3_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2630\,
            in2 => \_gnd_net_\,
            in3 => \N__2321\,
            lcout => \pwm_ctrZ0Z_3\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_2,
            carryout => pwm_ctr_cry_3,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_4_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2609\,
            in2 => \_gnd_net_\,
            in3 => \N__2318\,
            lcout => \pwm_ctrZ0Z_4\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_3,
            carryout => pwm_ctr_cry_4,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_5_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2582\,
            in2 => \_gnd_net_\,
            in3 => \N__2315\,
            lcout => \pwm_ctrZ0Z_5\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_4,
            carryout => pwm_ctr_cry_5,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_6_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2570\,
            in2 => \_gnd_net_\,
            in3 => \N__2312\,
            lcout => \pwm_ctrZ0Z_6\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_5,
            carryout => pwm_ctr_cry_6,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_7_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2558\,
            in2 => \_gnd_net_\,
            in3 => \N__2309\,
            lcout => \pwm_ctrZ0Z_7\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_6,
            carryout => pwm_ctr_cry_7,
            clk => \N__3217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_8_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2537\,
            in2 => \_gnd_net_\,
            in3 => \N__2306\,
            lcout => \pwm_ctrZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => pwm_ctr_cry_8,
            clk => \N__3216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_9_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2513\,
            in2 => \_gnd_net_\,
            in3 => \N__2342\,
            lcout => \pwm_ctrZ0Z_9\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_8,
            carryout => pwm_ctr_cry_9,
            clk => \N__3216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_10_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2501\,
            in2 => \_gnd_net_\,
            in3 => \N__2339\,
            lcout => \pwm_ctrZ0Z_10\,
            ltout => OPEN,
            carryin => pwm_ctr_cry_9,
            carryout => pwm_ctr_cry_10,
            clk => \N__3216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctr_11_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2489\,
            in2 => \_gnd_net_\,
            in3 => \N__2336\,
            lcout => \pwm_ctrZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIVDLC1_27_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000011011"
        )
    port map (
            in0 => \N__4410\,
            in1 => \N__3973\,
            in2 => \N__4533\,
            in3 => \N__4150\,
            lcout => pwm_g_1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNITBLC1_26_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110110001"
        )
    port map (
            in0 => \N__4149\,
            in1 => \N__3722\,
            in2 => \N__3811\,
            in3 => \N__4412\,
            lcout => pwm_g_1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNILGG11_29_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__4411\,
            in1 => \N__4151\,
            in2 => \_gnd_net_\,
            in3 => \N__3974\,
            lcout => pwm_g_1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_1_c_RNO_0_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000011011"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__2657\,
            in2 => \N__2474\,
            in3 => \N__2645\,
            lcout => OPEN,
            ltout => \N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_1_c_RNO_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4425\,
            in1 => \N__4162\,
            in2 => \N__2333\,
            in3 => \N__3614\,
            lcout => pwm_r_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIN5LC1_23_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000011011"
        )
    port map (
            in0 => \N__4426\,
            in1 => \N__4599\,
            in2 => \N__3493\,
            in3 => \N__4163\,
            lcout => pwm_g_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNI7D9M_21_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4836\,
            in2 => \N__3606\,
            in3 => \_gnd_net_\,
            lcout => \ctr_RNI7D9MZ0Z_21\,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => un34_r_val_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_1_c_RNIK0DV_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3595\,
            in2 => \N__4771\,
            in3 => \N__2366\,
            lcout => \un34_r_val_0_cry_1_c_RNIK0DVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_1,
            carryout => un34_r_val_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_2_c_RNIN4EV_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4758\,
            in2 => \N__3478\,
            in3 => \N__2363\,
            lcout => \un34_r_val_0_cry_2_c_RNIN4EVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_2,
            carryout => un34_r_val_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_3_c_RNIQ8FV_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3463\,
            in2 => \N__4721\,
            in3 => \N__2360\,
            lcout => \un34_r_val_0_cry_3_c_RNIQ8FVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_3,
            carryout => un34_r_val_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_4_c_RNITCGV_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4702\,
            in2 => \N__4600\,
            in3 => \N__2357\,
            lcout => \un34_r_val_0_cry_4_c_RNITCGVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_4,
            carryout => un34_r_val_0_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_5_c_RNI0HHV_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4588\,
            in2 => \N__3804\,
            in3 => \N__2354\,
            lcout => \un34_r_val_0_cry_5_c_RNI0HHVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_5,
            carryout => un34_r_val_0_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_6_c_RNI3LIV_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3789\,
            in2 => \N__4540\,
            in3 => \N__2351\,
            lcout => \un34_r_val_0_cry_6_c_RNI3LIVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_6,
            carryout => un34_r_val_0_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_7_c_RNI6PJV_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4532\,
            in2 => \N__3737\,
            in3 => \N__2348\,
            lcout => \un34_r_val_0_cry_7_c_RNI6PJVZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_7,
            carryout => un34_r_val_0_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_8_c_RNI9TKV_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3952\,
            in2 => \N__3723\,
            in3 => \N__2345\,
            lcout => \un34_r_val_0_cry_8_c_RNI9TKVZ0\,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => un34_r_val_0_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_9_c_RNIV0HK_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3972\,
            in3 => \N__2381\,
            lcout => \un34_r_val_0_cry_9_c_RNIV0HKZ0\,
            ltout => OPEN,
            carryin => un34_r_val_0_cry_9,
            carryout => un34_r_val_0_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un34_r_val_0_cry_10_THRU_LUT4_0_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2378\,
            lcout => \un34_r_val_0_cry_10_THRU_CO\,
            ltout => \un34_r_val_0_cry_10_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_11_c_RNO_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__3956\,
            in1 => \N__4376\,
            in2 => \N__2375\,
            in3 => \N__4096\,
            lcout => pwm_b_1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_5_c_RNO_0_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__3472\,
            in1 => \N__3420\,
            in2 => \N__4152\,
            in3 => \N__2819\,
            lcout => OPEN,
            ltout => \N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_5_c_RNO_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4362\,
            in1 => \N__4095\,
            in2 => \N__2372\,
            in3 => \N__4583\,
            lcout => pwm_r_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_3_c_RNO_0_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4090\,
            in1 => \N__3599\,
            in2 => \_gnd_net_\,
            in3 => \N__3555\,
            lcout => OPEN,
            ltout => \N_66_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_3_c_RNO_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4361\,
            in1 => \N__4091\,
            in2 => \N__2369\,
            in3 => \N__3473\,
            lcout => pwm_b_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIO5KC1_19_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000011101"
        )
    port map (
            in0 => \N__4064\,
            in1 => \N__2465\,
            in2 => \N__4413\,
            in3 => \N__3597\,
            lcout => pwm_g_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIM3KC1_18_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000011101"
        )
    port map (
            in0 => \N__4850\,
            in1 => \N__4349\,
            in2 => \N__4939\,
            in3 => \N__4066\,
            lcout => pwm_g_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_0_c_RNO_0_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__4062\,
            in1 => \N__4931\,
            in2 => \_gnd_net_\,
            in3 => \N__4847\,
            lcout => OPEN,
            ltout => \N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_0_c_RNO_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__4849\,
            in1 => \N__4348\,
            in2 => \N__2477\,
            in3 => \N__4065\,
            lcout => pwm_r_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIHVKC1_22_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101111010001"
        )
    port map (
            in0 => \N__4067\,
            in1 => \N__4769\,
            in2 => \N__4414\,
            in3 => \N__4851\,
            lcout => pwm_g_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIJ1LC1_21_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000110001011"
        )
    port map (
            in0 => \N__3598\,
            in1 => \N__4069\,
            in2 => \N__3488\,
            in3 => \N__4357\,
            lcout => pwm_g_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_1_c_RNO_0_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110011001"
        )
    port map (
            in0 => \N__4063\,
            in1 => \N__3596\,
            in2 => \_gnd_net_\,
            in3 => \N__4848\,
            lcout => OPEN,
            ltout => \un40_b_val_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_1_c_RNO_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010111000"
        )
    port map (
            in0 => \N__2466\,
            in1 => \N__4353\,
            in2 => \N__2444\,
            in3 => \N__4068\,
            lcout => pwm_b_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_0_c_inv_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3141\,
            in2 => \N__2441\,
            in3 => \N__2431\,
            lcout => pwm_ctr_i_0,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => pwm_g_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_1_c_inv_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2419\,
            in1 => \N__2408\,
            in2 => \N__3121\,
            in3 => \_gnd_net_\,
            lcout => pwm_ctr_i_1,
            ltout => OPEN,
            carryin => pwm_g_1_cry_0,
            carryout => pwm_g_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_2_c_inv_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2401\,
            in1 => \N__3075\,
            in2 => \N__2390\,
            in3 => \_gnd_net_\,
            lcout => pwm_ctr_i_2,
            ltout => OPEN,
            carryin => pwm_g_1_cry_1,
            carryout => pwm_g_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_3_c_inv_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2629\,
            in1 => \N__3042\,
            in2 => \N__2618\,
            in3 => \_gnd_net_\,
            lcout => pwm_ctr_i_3,
            ltout => OPEN,
            carryin => pwm_g_1_cry_2,
            carryout => pwm_g_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_4_c_inv_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3015\,
            in2 => \N__4664\,
            in3 => \N__2608\,
            lcout => pwm_ctr_i_4,
            ltout => OPEN,
            carryin => pwm_g_1_cry_3,
            carryout => pwm_g_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_5_c_inv_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2991\,
            in2 => \N__2597\,
            in3 => \N__2581\,
            lcout => pwm_ctr_i_5,
            ltout => OPEN,
            carryin => pwm_g_1_cry_4,
            carryout => pwm_g_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_6_c_inv_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3905\,
            in2 => \N__2973\,
            in3 => \N__2569\,
            lcout => pwm_ctr_i_6,
            ltout => OPEN,
            carryin => pwm_g_1_cry_5,
            carryout => pwm_g_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_7_c_inv_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2931\,
            in2 => \N__4649\,
            in3 => \N__2557\,
            lcout => pwm_ctr_i_7,
            ltout => OPEN,
            carryin => pwm_g_1_cry_6,
            carryout => pwm_g_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_8_c_inv_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3351\,
            in2 => \N__2546\,
            in3 => \N__2536\,
            lcout => pwm_ctr_i_8,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => pwm_g_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_9_c_inv_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3327\,
            in2 => \N__2525\,
            in3 => \N__2512\,
            lcout => pwm_ctr_i_9,
            ltout => OPEN,
            carryin => pwm_g_1_cry_8,
            carryout => pwm_g_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_10_c_inv_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2500\,
            in1 => \N__3288\,
            in2 => \N__2666\,
            in3 => \_gnd_net_\,
            lcout => pwm_ctr_i_10,
            ltout => OPEN,
            carryin => pwm_g_1_cry_9,
            carryout => pwm_g_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_1_cry_11_c_inv_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2488\,
            in1 => \N__3252\,
            in2 => \N__2693\,
            in3 => \_gnd_net_\,
            lcout => pwm_ctr_i_11,
            ltout => OPEN,
            carryin => pwm_g_1_cry_10,
            carryout => pwm_g_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_g_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2681\,
            lcout => \pwm_gZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_8_c_RNO_0_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4144\,
            in1 => \N__3803\,
            in2 => \_gnd_net_\,
            in3 => \N__3893\,
            lcout => OPEN,
            ltout => \N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_8_c_RNO_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4423\,
            in1 => \N__3730\,
            in2 => \N__2669\,
            in3 => \N__4145\,
            lcout => pwm_b_1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIKFG11_28_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__3731\,
            in1 => \_gnd_net_\,
            in2 => \N__4224\,
            in3 => \N__4424\,
            lcout => pwm_g_1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_0_c_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4865\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => un33_r_val_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_0_THRU_LUT4_0_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2656\,
            in2 => \N__2773\,
            in3 => \N__2639\,
            lcout => \un33_r_val_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_0,
            carryout => un33_r_val_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_1_THRU_LUT4_0_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2755\,
            in2 => \N__4899\,
            in3 => \N__2636\,
            lcout => \un33_r_val_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_1,
            carryout => un33_r_val_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_2_THRU_LUT4_0_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2758\,
            in2 => \N__3556\,
            in3 => \N__2633\,
            lcout => \un33_r_val_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_2,
            carryout => un33_r_val_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_3_THRU_LUT4_0_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2756\,
            in2 => \N__3652\,
            in3 => \N__2822\,
            lcout => \un33_r_val_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_3,
            carryout => un33_r_val_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_4_THRU_LUT4_0_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2759\,
            in2 => \N__3424\,
            in3 => \N__2810\,
            lcout => \un33_r_val_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_4,
            carryout => un33_r_val_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_5_THRU_LUT4_0_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2757\,
            in2 => \N__3840\,
            in3 => \N__2807\,
            lcout => \un33_r_val_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_5,
            carryout => un33_r_val_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_6_THRU_LUT4_0_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2760\,
            in2 => \N__4629\,
            in3 => \N__2804\,
            lcout => \un33_r_val_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_6,
            carryout => un33_r_val_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_7_THRU_LUT4_0_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2761\,
            in2 => \N__3882\,
            in3 => \N__2801\,
            lcout => \un33_r_val_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => un33_r_val_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_8_THRU_LUT4_0_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2762\,
            in2 => \N__3190\,
            in3 => \N__2711\,
            lcout => \un33_r_val_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => un33_r_val_cry_8,
            carryout => un33_r_val_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_10_c_RNO_0_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2879\,
            in3 => \N__2708\,
            lcout => \pwm_r_1_cry_10_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => un33_r_val_cry_9,
            carryout => un33_r_val_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un33_r_val_cry_10_THRU_LUT4_0_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2705\,
            lcout => OPEN,
            ltout => \un33_r_val_cry_10_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_11_c_RNO_0_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2702\,
            in3 => \N__2699\,
            lcout => \pwm_r_1_cry_11_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_4_c_RNO_0_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__4793\,
            in1 => \N__3648\,
            in2 => \N__4258\,
            in3 => \N__2864\,
            lcout => OPEN,
            ltout => \N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_4_c_RNO_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4458\,
            in1 => \N__4221\,
            in2 => \N__2858\,
            in3 => \N__4726\,
            lcout => pwm_r_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_0_c_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2855\,
            in2 => \N__3149\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_27_0_\,
            carryout => pwm_r_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_1_c_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2849\,
            in2 => \N__3122\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_0,
            carryout => pwm_r_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_2_c_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3083\,
            in2 => \N__3626\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_1,
            carryout => pwm_r_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_3_c_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3050\,
            in2 => \N__3524\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_2,
            carryout => pwm_r_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_4_c_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3026\,
            in2 => \N__2840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_3,
            carryout => pwm_r_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_5_c_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2999\,
            in2 => \N__2831\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_4,
            carryout => pwm_r_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_6_c_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2975\,
            in2 => \N__3503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_5,
            carryout => pwm_r_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_7_c_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2945\,
            in2 => \N__3374\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_6,
            carryout => pwm_r_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_8_c_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3359\,
            in2 => \N__3854\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_28_0_\,
            carryout => pwm_r_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_9_c_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3335\,
            in2 => \N__2888\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_8,
            carryout => pwm_r_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_10_c_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3662\,
            in2 => \N__3302\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_9,
            carryout => pwm_r_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_11_c_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3262\,
            in2 => \N__3914\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_r_1_cry_10,
            carryout => pwm_r_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2915\,
            lcout => \pwm_rZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_9_c_RNO_0_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__4528\,
            in1 => \N__3186\,
            in2 => \N__4226\,
            in3 => \N__2900\,
            lcout => OPEN,
            ltout => \N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_9_c_RNO_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4419\,
            in1 => \N__4159\,
            in2 => \N__2891\,
            in3 => \N__3981\,
            lcout => pwm_r_1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_10_c_RNO_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__3724\,
            in1 => \N__4418\,
            in2 => \N__4225\,
            in3 => \N__2878\,
            lcout => pwm_b_1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_0_c_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4913\,
            in2 => \N__3148\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => pwm_b_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_1_c_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3111\,
            in2 => \N__3092\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_0,
            carryout => pwm_b_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_2_c_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4802\,
            in2 => \N__3082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_1,
            carryout => pwm_b_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_3_c_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3059\,
            in2 => \N__3049\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_2,
            carryout => pwm_b_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_4_c_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4949\,
            in2 => \N__3022\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_3,
            carryout => pwm_b_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_5_c_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3398\,
            in2 => \N__2998\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_4,
            carryout => pwm_b_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_6_c_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3746\,
            in2 => \N__2974\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_5,
            carryout => pwm_b_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_7_c_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3992\,
            in2 => \N__2944\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_6,
            carryout => pwm_b_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_8_c_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3365\,
            in2 => \N__3358\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_30_0_\,
            carryout => pwm_b_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_9_c_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3164\,
            in2 => \N__3334\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_8,
            carryout => pwm_b_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_10_c_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3311\,
            in2 => \N__3301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_9,
            carryout => pwm_b_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_11_c_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3272\,
            in2 => \N__3263\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => pwm_b_1_cry_10,
            carryout => pwm_b_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3236\,
            lcout => \pwm_bZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_9_c_RNO_0_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4222\,
            in1 => \N__4539\,
            in2 => \_gnd_net_\,
            in3 => \N__3194\,
            lcout => OPEN,
            ltout => \N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_9_c_RNO_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4459\,
            in1 => \N__4223\,
            in2 => \N__3167\,
            in3 => \N__3985\,
            lcout => pwm_b_1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_2_c_RNO_0_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000011101"
        )
    port map (
            in0 => \N__4906\,
            in1 => \N__4205\,
            in2 => \N__4873\,
            in3 => \N__3158\,
            lcout => OPEN,
            ltout => \N_89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_2_c_RNO_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4434\,
            in1 => \N__4217\,
            in2 => \N__3152\,
            in3 => \N__4796\,
            lcout => pwm_r_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_3_c_RNO_0_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__3613\,
            in1 => \N__3560\,
            in2 => \N__4254\,
            in3 => \N__3533\,
            lcout => OPEN,
            ltout => \N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_3_c_RNO_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__3494\,
            in1 => \N__4435\,
            in2 => \N__3527\,
            in3 => \N__4209\,
            lcout => pwm_r_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_6_c_RNO_0_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__4724\,
            in1 => \N__3841\,
            in2 => \N__4259\,
            in3 => \N__3512\,
            lcout => OPEN,
            ltout => \N_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_6_c_RNO_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__3812\,
            in1 => \N__4233\,
            in2 => \N__3506\,
            in3 => \N__4461\,
            lcout => pwm_r_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_5_c_RNO_0_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__3489\,
            in2 => \_gnd_net_\,
            in3 => \N__3425\,
            lcout => OPEN,
            ltout => \N_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_5_c_RNO_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__4603\,
            in1 => \N__4460\,
            in2 => \N__3401\,
            in3 => \N__4228\,
            lcout => pwm_b_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_7_c_RNO_0_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001000100111"
        )
    port map (
            in0 => \N__4232\,
            in1 => \N__4604\,
            in2 => \N__3386\,
            in3 => \N__4633\,
            lcout => OPEN,
            ltout => \N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_7_c_RNO_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__4541\,
            in1 => \N__4234\,
            in2 => \N__3377\,
            in3 => \N__4462\,
            lcout => pwm_r_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_11_c_RNO_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000010"
        )
    port map (
            in0 => \N__4253\,
            in1 => \N__4442\,
            in2 => \N__3986\,
            in3 => \N__3920\,
            lcout => pwm_r_1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIP7LC1_24_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000011011"
        )
    port map (
            in0 => \N__4723\,
            in1 => \N__4244\,
            in2 => \N__4463\,
            in3 => \N__3805\,
            lcout => pwm_g_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_8_c_RNO_0_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010011"
        )
    port map (
            in0 => \N__3807\,
            in1 => \N__3889\,
            in2 => \N__4261\,
            in3 => \N__3863\,
            lcout => OPEN,
            ltout => \N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_8_c_RNO_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__4440\,
            in1 => \N__4249\,
            in2 => \N__3857\,
            in3 => \N__3735\,
            lcout => pwm_r_1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_6_c_RNO_0_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4243\,
            in1 => \N__4722\,
            in2 => \_gnd_net_\,
            in3 => \N__3845\,
            lcout => OPEN,
            ltout => \N_69_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_6_c_RNO_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4439\,
            in1 => \N__4245\,
            in2 => \N__3815\,
            in3 => \N__3806\,
            lcout => pwm_b_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_r_1_cry_10_c_RNO_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__3736\,
            in1 => \N__4441\,
            in2 => \N__4262\,
            in3 => \N__3668\,
            lcout => pwm_r_1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_4_c_RNO_0_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__4255\,
            in1 => \N__4784\,
            in2 => \_gnd_net_\,
            in3 => \N__3656\,
            lcout => OPEN,
            ltout => \N_67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_4_c_RNO_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4465\,
            in1 => \N__4257\,
            in2 => \N__3629\,
            in3 => \N__4725\,
            lcout => pwm_b_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_0_c_RNO_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001101"
        )
    port map (
            in0 => \N__4464\,
            in1 => \N__4943\,
            in2 => \N__4877\,
            in3 => \N__4256\,
            lcout => pwm_b_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_2_c_RNO_0_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__4235\,
            in1 => \N__4907\,
            in2 => \_gnd_net_\,
            in3 => \N__4872\,
            lcout => OPEN,
            ltout => \N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_2_c_RNO_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__4471\,
            in1 => \N__4239\,
            in2 => \N__4805\,
            in3 => \N__4794\,
            lcout => pwm_b_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIL3LC1_22_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000100111"
        )
    port map (
            in0 => \N__4795\,
            in1 => \N__4470\,
            in2 => \N__4260\,
            in3 => \N__4727\,
            lcout => pwm_g_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ctr_RNIR9LC1_25_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101111010001"
        )
    port map (
            in0 => \N__4240\,
            in1 => \N__4534\,
            in2 => \N__4472\,
            in3 => \N__4602\,
            lcout => pwm_g_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_7_c_RNO_0_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__4241\,
            in1 => \N__4634\,
            in2 => \_gnd_net_\,
            in3 => \N__4601\,
            lcout => OPEN,
            ltout => \N_70_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_b_1_cry_7_c_RNO_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__4535\,
            in1 => \N__4469\,
            in2 => \N__4265\,
            in3 => \N__4242\,
            lcout => pwm_b_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
