// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 6 2018 12:49:44

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    RGB2,
    RGB1,
    RGB0);

    output RGB2;
    output RGB1;
    output RGB0;

    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4939;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4920;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4885;
    wire N__4882;
    wire N__4877;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4852;
    wire N__4851;
    wire N__4850;
    wire N__4849;
    wire N__4848;
    wire N__4847;
    wire N__4844;
    wire N__4837;
    wire N__4836;
    wire N__4833;
    wire N__4822;
    wire N__4817;
    wire N__4814;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4793;
    wire N__4790;
    wire N__4785;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4771;
    wire N__4770;
    wire N__4769;
    wire N__4766;
    wire N__4759;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4738;
    wire N__4727;
    wire N__4726;
    wire N__4725;
    wire N__4724;
    wire N__4723;
    wire N__4722;
    wire N__4721;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4703;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4684;
    wire N__4679;
    wire N__4672;
    wire N__4669;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4633;
    wire N__4630;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4604;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4599;
    wire N__4594;
    wire N__4589;
    wire N__4588;
    wire N__4585;
    wire N__4584;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4552;
    wire N__4541;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4535;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4509;
    wire N__4508;
    wire N__4505;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4484;
    wire N__4479;
    wire N__4472;
    wire N__4471;
    wire N__4470;
    wire N__4469;
    wire N__4466;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4460;
    wire N__4459;
    wire N__4458;
    wire N__4453;
    wire N__4448;
    wire N__4443;
    wire N__4442;
    wire N__4441;
    wire N__4440;
    wire N__4439;
    wire N__4436;
    wire N__4435;
    wire N__4434;
    wire N__4427;
    wire N__4426;
    wire N__4425;
    wire N__4424;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4418;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4411;
    wire N__4410;
    wire N__4407;
    wire N__4402;
    wire N__4391;
    wire N__4386;
    wire N__4383;
    wire N__4378;
    wire N__4377;
    wire N__4376;
    wire N__4371;
    wire N__4368;
    wire N__4363;
    wire N__4362;
    wire N__4361;
    wire N__4358;
    wire N__4357;
    wire N__4354;
    wire N__4353;
    wire N__4350;
    wire N__4349;
    wire N__4348;
    wire N__4341;
    wire N__4334;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4313;
    wire N__4308;
    wire N__4305;
    wire N__4292;
    wire N__4287;
    wire N__4284;
    wire N__4265;
    wire N__4262;
    wire N__4261;
    wire N__4260;
    wire N__4259;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4249;
    wire N__4246;
    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4236;
    wire N__4235;
    wire N__4234;
    wire N__4233;
    wire N__4232;
    wire N__4229;
    wire N__4228;
    wire N__4227;
    wire N__4226;
    wire N__4225;
    wire N__4224;
    wire N__4223;
    wire N__4222;
    wire N__4221;
    wire N__4218;
    wire N__4217;
    wire N__4210;
    wire N__4209;
    wire N__4206;
    wire N__4205;
    wire N__4190;
    wire N__4177;
    wire N__4164;
    wire N__4163;
    wire N__4162;
    wire N__4161;
    wire N__4160;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4152;
    wire N__4151;
    wire N__4150;
    wire N__4149;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4139;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4121;
    wire N__4114;
    wire N__4107;
    wire N__4104;
    wire N__4097;
    wire N__4096;
    wire N__4095;
    wire N__4092;
    wire N__4091;
    wire N__4090;
    wire N__4083;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4064;
    wire N__4063;
    wire N__4062;
    wire N__4059;
    wire N__4050;
    wire N__4045;
    wire N__4034;
    wire N__4025;
    wire N__4008;
    wire N__4003;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3985;
    wire N__3982;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3974;
    wire N__3973;
    wire N__3972;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3957;
    wire N__3956;
    wire N__3953;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3938;
    wire N__3931;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3882;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3841;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3815;
    wire N__3812;
    wire N__3811;
    wire N__3808;
    wire N__3807;
    wire N__3806;
    wire N__3805;
    wire N__3804;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3790;
    wire N__3789;
    wire N__3786;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3774;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3758;
    wire N__3755;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3736;
    wire N__3735;
    wire N__3732;
    wire N__3731;
    wire N__3730;
    wire N__3725;
    wire N__3724;
    wire N__3723;
    wire N__3722;
    wire N__3719;
    wire N__3718;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3687;
    wire N__3684;
    wire N__3679;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3652;
    wire N__3649;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3606;
    wire N__3605;
    wire N__3600;
    wire N__3599;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3576;
    wire N__3571;
    wire N__3560;
    wire N__3557;
    wire N__3556;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3512;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3489;
    wire N__3488;
    wire N__3485;
    wire N__3482;
    wire N__3479;
    wire N__3478;
    wire N__3477;
    wire N__3474;
    wire N__3473;
    wire N__3472;
    wire N__3469;
    wire N__3464;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3438;
    wire N__3425;
    wire N__3424;
    wire N__3421;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3335;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3223;
    wire N__3222;
    wire N__3221;
    wire N__3220;
    wire N__3219;
    wire N__3218;
    wire N__3217;
    wire N__3216;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3190;
    wire N__3187;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3149;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3122;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3097;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3026;
    wire N__3023;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__2999;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2975;
    wire N__2974;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2945;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2878;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2813;
    wire N__2810;
    wire N__2807;
    wire N__2804;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2794;
    wire N__2791;
    wire N__2790;
    wire N__2787;
    wire N__2786;
    wire N__2783;
    wire N__2780;
    wire N__2777;
    wire N__2774;
    wire N__2773;
    wire N__2770;
    wire N__2763;
    wire N__2762;
    wire N__2761;
    wire N__2760;
    wire N__2759;
    wire N__2758;
    wire N__2757;
    wire N__2756;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2733;
    wire N__2724;
    wire N__2711;
    wire N__2708;
    wire N__2705;
    wire N__2702;
    wire N__2699;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2678;
    wire N__2675;
    wire N__2672;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2657;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2645;
    wire N__2642;
    wire N__2639;
    wire N__2636;
    wire N__2633;
    wire N__2630;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2618;
    wire N__2615;
    wire N__2612;
    wire N__2609;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2597;
    wire N__2594;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2570;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2558;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2546;
    wire N__2543;
    wire N__2540;
    wire N__2537;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2501;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2489;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2468;
    wire N__2467;
    wire N__2466;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2454;
    wire N__2451;
    wire N__2444;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2420;
    wire N__2419;
    wire N__2416;
    wire N__2413;
    wire N__2408;
    wire N__2405;
    wire N__2402;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2378;
    wire N__2375;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2360;
    wire N__2357;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2270;
    wire N__2267;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2240;
    wire N__2237;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2225;
    wire N__2222;
    wire N__2219;
    wire N__2216;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2183;
    wire N__2180;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2168;
    wire N__2165;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire N__2150;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2114;
    wire N__2111;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire VCCG0;
    wire GNDG0;
    wire ctrZ0Z_0;
    wire bfn_1_25_0_;
    wire ctrZ0Z_1;
    wire ctr_cry_0;
    wire ctrZ0Z_2;
    wire ctr_cry_1;
    wire ctrZ0Z_3;
    wire ctr_cry_2;
    wire ctrZ0Z_4;
    wire ctr_cry_3;
    wire ctrZ0Z_5;
    wire ctr_cry_4;
    wire ctrZ0Z_6;
    wire ctr_cry_5;
    wire ctrZ0Z_7;
    wire ctr_cry_6;
    wire ctr_cry_7;
    wire ctrZ0Z_8;
    wire bfn_1_26_0_;
    wire ctrZ0Z_9;
    wire ctr_cry_8;
    wire ctrZ0Z_10;
    wire ctr_cry_9;
    wire ctrZ0Z_11;
    wire ctr_cry_10;
    wire ctrZ0Z_12;
    wire ctr_cry_11;
    wire ctrZ0Z_13;
    wire ctr_cry_12;
    wire ctrZ0Z_14;
    wire ctr_cry_13;
    wire ctrZ0Z_15;
    wire ctr_cry_14;
    wire ctr_cry_15;
    wire ctrZ0Z_16;
    wire bfn_1_27_0_;
    wire ctrZ0Z_17;
    wire ctr_cry_16;
    wire ctr_cry_17;
    wire ctr_cry_18;
    wire ctr_cry_19;
    wire ctr_cry_20;
    wire ctr_cry_21;
    wire ctr_cry_22;
    wire ctr_cry_23;
    wire bfn_1_28_0_;
    wire ctr_cry_24;
    wire ctr_cry_25;
    wire ctr_cry_26;
    wire ctr_cry_27;
    wire ctr_cry_28;
    wire ctr_cry_29;
    wire ctr_cry_30;
    wire bfn_1_29_0_;
    wire pwm_ctr_cry_0;
    wire pwm_ctr_cry_1;
    wire pwm_ctr_cry_2;
    wire pwm_ctr_cry_3;
    wire pwm_ctr_cry_4;
    wire pwm_ctr_cry_5;
    wire pwm_ctr_cry_6;
    wire pwm_ctr_cry_7;
    wire bfn_1_30_0_;
    wire pwm_ctr_cry_8;
    wire pwm_ctr_cry_9;
    wire pwm_ctr_cry_10;
    wire N_88_cascade_;
    wire bfn_2_26_0_;
    wire un34_r_val_0_cry_1;
    wire un34_r_val_0_cry_2;
    wire un34_r_val_0_cry_3;
    wire un34_r_val_0_cry_4;
    wire un34_r_val_0_cry_5;
    wire un34_r_val_0_cry_6;
    wire un34_r_val_0_cry_7;
    wire un34_r_val_0_cry_8;
    wire bfn_2_27_0_;
    wire un34_r_val_0_cry_9;
    wire un34_r_val_0_cry_10;
    wire un34_r_val_0_cry_10_THRU_CO_cascade_;
    wire N_92_cascade_;
    wire N_66_cascade_;
    wire N_87_cascade_;
    wire ctrZ0Z_19;
    wire un40_b_val_3_ns_1_1_cascade_;
    wire pwm_g_1_0;
    wire pwm_ctrZ0Z_0;
    wire bfn_2_29_0_;
    wire pwm_ctrZ0Z_1;
    wire pwm_g_1_1;
    wire pwm_g_1_cry_0;
    wire pwm_ctrZ0Z_2;
    wire pwm_g_1_2;
    wire pwm_g_1_cry_1;
    wire pwm_ctrZ0Z_3;
    wire pwm_g_1_3;
    wire pwm_g_1_cry_2;
    wire pwm_ctrZ0Z_4;
    wire pwm_g_1_cry_3;
    wire pwm_g_1_5;
    wire pwm_ctrZ0Z_5;
    wire pwm_g_1_cry_4;
    wire pwm_ctrZ0Z_6;
    wire pwm_g_1_cry_5;
    wire pwm_ctrZ0Z_7;
    wire pwm_g_1_cry_6;
    wire pwm_g_1_cry_7;
    wire pwm_g_1_8;
    wire pwm_ctrZ0Z_8;
    wire bfn_2_30_0_;
    wire pwm_g_1_9;
    wire pwm_ctrZ0Z_9;
    wire pwm_g_1_cry_8;
    wire pwm_ctrZ0Z_10;
    wire pwm_g_1_cry_9;
    wire pwm_ctrZ0Z_11;
    wire pwm_g_1_11;
    wire pwm_g_1_cry_10;
    wire pwm_g_1;
    wire pwm_gZ0;
    wire N_71_cascade_;
    wire pwm_g_1_10;
    wire bfn_3_25_0_;
    wire ctr_RNI7D9MZ0Z_21;
    wire un33_r_val_cry_0_THRU_CO;
    wire un33_r_val_cry_0;
    wire un33_r_val_cry_1;
    wire un33_r_val_cry_2;
    wire un33_r_val_cry_3;
    wire un33_r_val_cry_4_THRU_CO;
    wire un33_r_val_cry_4;
    wire un33_r_val_cry_5;
    wire un33_r_val_cry_6;
    wire un33_r_val_cry_7;
    wire bfn_3_26_0_;
    wire CONSTANT_ONE_NET;
    wire un33_r_val_cry_8;
    wire un33_r_val_cry_9;
    wire un33_r_val_cry_10;
    wire un33_r_val_cry_10_THRU_CO_cascade_;
    wire un34_r_val_0_cry_10_THRU_CO;
    wire un33_r_val_cry_3_THRU_CO;
    wire N_91_cascade_;
    wire pwm_r_1_0;
    wire bfn_3_27_0_;
    wire pwm_r_1_1;
    wire pwm_r_1_cry_0;
    wire pwm_r_1_cry_1;
    wire pwm_r_1_cry_2;
    wire pwm_r_1_4;
    wire pwm_r_1_cry_3;
    wire pwm_r_1_5;
    wire pwm_r_1_cry_4;
    wire pwm_r_1_cry_5;
    wire pwm_r_1_cry_6;
    wire pwm_r_1_cry_7;
    wire bfn_3_28_0_;
    wire pwm_r_1_cry_8;
    wire pwm_r_1_cry_9;
    wire pwm_r_1_cry_10;
    wire pwm_r_1;
    wire pwm_rZ0;
    wire un33_r_val_cry_8_THRU_CO;
    wire N_96_cascade_;
    wire pwm_r_1_9;
    wire un34_r_val_0_cry_9_c_RNIV0HKZ0;
    wire pwm_ctr_i_0;
    wire bfn_3_29_0_;
    wire pwm_ctr_i_1;
    wire pwm_b_1_1;
    wire pwm_b_1_cry_0;
    wire pwm_ctr_i_2;
    wire pwm_b_1_cry_1;
    wire pwm_b_1_3;
    wire pwm_ctr_i_3;
    wire pwm_b_1_cry_2;
    wire pwm_ctr_i_4;
    wire pwm_b_1_cry_3;
    wire pwm_ctr_i_5;
    wire pwm_b_1_cry_4;
    wire pwm_ctr_i_6;
    wire pwm_b_1_cry_5;
    wire pwm_ctr_i_7;
    wire pwm_b_1_cry_6;
    wire pwm_b_1_cry_7;
    wire pwm_b_1_8;
    wire pwm_ctr_i_8;
    wire bfn_3_30_0_;
    wire pwm_ctr_i_9;
    wire pwm_b_1_cry_8;
    wire pwm_b_1_10;
    wire pwm_ctr_i_10;
    wire pwm_b_1_cry_9;
    wire pwm_b_1_11;
    wire pwm_ctr_i_11;
    wire pwm_b_1_cry_10;
    wire pwm_b_1;
    wire pwm_bZ0;
    wire clk;
    wire un34_r_val_0_cry_8_c_RNI9TKVZ0;
    wire N_72_cascade_;
    wire pwm_b_1_9;
    wire un33_r_val_cry_1_THRU_CO;
    wire N_89_cascade_;
    wire pwm_r_1_2;
    wire ctrZ0Z_21;
    wire un34_r_val_0_cry_2_c_RNIN4EVZ0;
    wire un33_r_val_cry_2_THRU_CO;
    wire N_90_cascade_;
    wire pwm_r_1_3;
    wire un33_r_val_cry_5_THRU_CO;
    wire N_93_cascade_;
    wire pwm_r_1_6;
    wire ctrZ0Z_23;
    wire un34_r_val_0_cry_4_c_RNITCGVZ0;
    wire N_68_cascade_;
    wire pwm_b_1_5;
    wire un33_r_val_cry_6_THRU_CO;
    wire N_94_cascade_;
    wire pwm_r_1_7;
    wire ctrZ0Z_29;
    wire pwm_r_1_cry_11_c_RNOZ0Z_0;
    wire pwm_r_1_11;
    wire pwm_g_1_6;
    wire un34_r_val_0_cry_7_c_RNI6PJVZ0;
    wire un33_r_val_cry_7_THRU_CO;
    wire N_95_cascade_;
    wire pwm_r_1_8;
    wire un34_r_val_0_cry_5_c_RNI0HHVZ0;
    wire N_69_cascade_;
    wire ctrZ0Z_26;
    wire pwm_b_1_6;
    wire ctrZ0Z_28;
    wire pwm_r_1_cry_10_c_RNOZ0Z_0;
    wire pwm_r_1_10;
    wire un34_r_val_0_cry_3_c_RNIQ8FVZ0;
    wire N_67_cascade_;
    wire pwm_b_1_4;
    wire ctrZ0Z_18;
    wire pwm_b_1_0;
    wire un34_r_val_0_cry_1_c_RNIK0DVZ0;
    wire ctrZ0Z_20;
    wire N_65_cascade_;
    wire pwm_b_1_2;
    wire ctrZ0Z_22;
    wire ctrZ0Z_24;
    wire pwm_g_1_4;
    wire pwm_g_1_7;
    wire un34_r_val_0_cry_6_c_RNI3LIVZ0;
    wire ctrZ0Z_25;
    wire ctrZ0Z_27;
    wire ctrZ0Z_31;
    wire N_70_cascade_;
    wire ctrZ0Z_30;
    wire pwm_b_1_7;
    wire _gnd_net_;

    InMux I__1133 (
            .O(N__4949),
            .I(N__4946));
    LocalMux I__1132 (
            .O(N__4946),
            .I(pwm_b_1_4));
    InMux I__1131 (
            .O(N__4943),
            .I(N__4940));
    LocalMux I__1130 (
            .O(N__4940),
            .I(N__4935));
    CascadeMux I__1129 (
            .O(N__4939),
            .I(N__4932));
    InMux I__1128 (
            .O(N__4938),
            .I(N__4928));
    Span4Mux_h I__1127 (
            .O(N__4935),
            .I(N__4925));
    InMux I__1126 (
            .O(N__4932),
            .I(N__4920));
    InMux I__1125 (
            .O(N__4931),
            .I(N__4920));
    LocalMux I__1124 (
            .O(N__4928),
            .I(ctrZ0Z_18));
    Odrv4 I__1123 (
            .O(N__4925),
            .I(ctrZ0Z_18));
    LocalMux I__1122 (
            .O(N__4920),
            .I(ctrZ0Z_18));
    InMux I__1121 (
            .O(N__4913),
            .I(N__4910));
    LocalMux I__1120 (
            .O(N__4910),
            .I(pwm_b_1_0));
    InMux I__1119 (
            .O(N__4907),
            .I(N__4903));
    InMux I__1118 (
            .O(N__4906),
            .I(N__4900));
    LocalMux I__1117 (
            .O(N__4903),
            .I(N__4896));
    LocalMux I__1116 (
            .O(N__4900),
            .I(N__4893));
    CascadeMux I__1115 (
            .O(N__4899),
            .I(N__4890));
    Span4Mux_v I__1114 (
            .O(N__4896),
            .I(N__4885));
    Span4Mux_v I__1113 (
            .O(N__4893),
            .I(N__4885));
    InMux I__1112 (
            .O(N__4890),
            .I(N__4882));
    Odrv4 I__1111 (
            .O(N__4885),
            .I(un34_r_val_0_cry_1_c_RNIK0DVZ0));
    LocalMux I__1110 (
            .O(N__4882),
            .I(un34_r_val_0_cry_1_c_RNIK0DVZ0));
    CascadeMux I__1109 (
            .O(N__4877),
            .I(N__4874));
    InMux I__1108 (
            .O(N__4874),
            .I(N__4869));
    CascadeMux I__1107 (
            .O(N__4873),
            .I(N__4866));
    InMux I__1106 (
            .O(N__4872),
            .I(N__4862));
    LocalMux I__1105 (
            .O(N__4869),
            .I(N__4859));
    InMux I__1104 (
            .O(N__4866),
            .I(N__4856));
    InMux I__1103 (
            .O(N__4865),
            .I(N__4853));
    LocalMux I__1102 (
            .O(N__4862),
            .I(N__4844));
    Span4Mux_v I__1101 (
            .O(N__4859),
            .I(N__4837));
    LocalMux I__1100 (
            .O(N__4856),
            .I(N__4837));
    LocalMux I__1099 (
            .O(N__4853),
            .I(N__4837));
    InMux I__1098 (
            .O(N__4852),
            .I(N__4833));
    InMux I__1097 (
            .O(N__4851),
            .I(N__4822));
    InMux I__1096 (
            .O(N__4850),
            .I(N__4822));
    InMux I__1095 (
            .O(N__4849),
            .I(N__4822));
    InMux I__1094 (
            .O(N__4848),
            .I(N__4822));
    InMux I__1093 (
            .O(N__4847),
            .I(N__4822));
    Span4Mux_h I__1092 (
            .O(N__4844),
            .I(N__4817));
    Span4Mux_h I__1091 (
            .O(N__4837),
            .I(N__4817));
    InMux I__1090 (
            .O(N__4836),
            .I(N__4814));
    LocalMux I__1089 (
            .O(N__4833),
            .I(ctrZ0Z_20));
    LocalMux I__1088 (
            .O(N__4822),
            .I(ctrZ0Z_20));
    Odrv4 I__1087 (
            .O(N__4817),
            .I(ctrZ0Z_20));
    LocalMux I__1086 (
            .O(N__4814),
            .I(ctrZ0Z_20));
    CascadeMux I__1085 (
            .O(N__4805),
            .I(N_65_cascade_));
    InMux I__1084 (
            .O(N__4802),
            .I(N__4799));
    LocalMux I__1083 (
            .O(N__4799),
            .I(pwm_b_1_2));
    InMux I__1082 (
            .O(N__4796),
            .I(N__4790));
    InMux I__1081 (
            .O(N__4795),
            .I(N__4785));
    InMux I__1080 (
            .O(N__4794),
            .I(N__4785));
    InMux I__1079 (
            .O(N__4793),
            .I(N__4781));
    LocalMux I__1078 (
            .O(N__4790),
            .I(N__4778));
    LocalMux I__1077 (
            .O(N__4785),
            .I(N__4775));
    InMux I__1076 (
            .O(N__4784),
            .I(N__4772));
    LocalMux I__1075 (
            .O(N__4781),
            .I(N__4766));
    Span4Mux_v I__1074 (
            .O(N__4778),
            .I(N__4759));
    Span4Mux_s2_v I__1073 (
            .O(N__4775),
            .I(N__4759));
    LocalMux I__1072 (
            .O(N__4772),
            .I(N__4759));
    CascadeMux I__1071 (
            .O(N__4771),
            .I(N__4755));
    InMux I__1070 (
            .O(N__4770),
            .I(N__4752));
    InMux I__1069 (
            .O(N__4769),
            .I(N__4749));
    Span4Mux_h I__1068 (
            .O(N__4766),
            .I(N__4746));
    Span4Mux_h I__1067 (
            .O(N__4759),
            .I(N__4743));
    InMux I__1066 (
            .O(N__4758),
            .I(N__4738));
    InMux I__1065 (
            .O(N__4755),
            .I(N__4738));
    LocalMux I__1064 (
            .O(N__4752),
            .I(ctrZ0Z_22));
    LocalMux I__1063 (
            .O(N__4749),
            .I(ctrZ0Z_22));
    Odrv4 I__1062 (
            .O(N__4746),
            .I(ctrZ0Z_22));
    Odrv4 I__1061 (
            .O(N__4743),
            .I(ctrZ0Z_22));
    LocalMux I__1060 (
            .O(N__4738),
            .I(ctrZ0Z_22));
    InMux I__1059 (
            .O(N__4727),
            .I(N__4717));
    InMux I__1058 (
            .O(N__4726),
            .I(N__4714));
    InMux I__1057 (
            .O(N__4725),
            .I(N__4711));
    InMux I__1056 (
            .O(N__4724),
            .I(N__4708));
    InMux I__1055 (
            .O(N__4723),
            .I(N__4703));
    InMux I__1054 (
            .O(N__4722),
            .I(N__4703));
    CascadeMux I__1053 (
            .O(N__4721),
            .I(N__4699));
    InMux I__1052 (
            .O(N__4720),
            .I(N__4696));
    LocalMux I__1051 (
            .O(N__4717),
            .I(N__4693));
    LocalMux I__1050 (
            .O(N__4714),
            .I(N__4684));
    LocalMux I__1049 (
            .O(N__4711),
            .I(N__4684));
    LocalMux I__1048 (
            .O(N__4708),
            .I(N__4684));
    LocalMux I__1047 (
            .O(N__4703),
            .I(N__4684));
    InMux I__1046 (
            .O(N__4702),
            .I(N__4679));
    InMux I__1045 (
            .O(N__4699),
            .I(N__4679));
    LocalMux I__1044 (
            .O(N__4696),
            .I(N__4672));
    Span4Mux_s2_v I__1043 (
            .O(N__4693),
            .I(N__4672));
    Span4Mux_v I__1042 (
            .O(N__4684),
            .I(N__4672));
    LocalMux I__1041 (
            .O(N__4679),
            .I(N__4669));
    Odrv4 I__1040 (
            .O(N__4672),
            .I(ctrZ0Z_24));
    Odrv4 I__1039 (
            .O(N__4669),
            .I(ctrZ0Z_24));
    CascadeMux I__1038 (
            .O(N__4664),
            .I(N__4661));
    InMux I__1037 (
            .O(N__4661),
            .I(N__4658));
    LocalMux I__1036 (
            .O(N__4658),
            .I(N__4655));
    Span4Mux_s3_h I__1035 (
            .O(N__4655),
            .I(N__4652));
    Odrv4 I__1034 (
            .O(N__4652),
            .I(pwm_g_1_4));
    CascadeMux I__1033 (
            .O(N__4649),
            .I(N__4646));
    InMux I__1032 (
            .O(N__4646),
            .I(N__4643));
    LocalMux I__1031 (
            .O(N__4643),
            .I(N__4640));
    Span4Mux_h I__1030 (
            .O(N__4640),
            .I(N__4637));
    Odrv4 I__1029 (
            .O(N__4637),
            .I(pwm_g_1_7));
    InMux I__1028 (
            .O(N__4634),
            .I(N__4630));
    InMux I__1027 (
            .O(N__4633),
            .I(N__4626));
    LocalMux I__1026 (
            .O(N__4630),
            .I(N__4623));
    CascadeMux I__1025 (
            .O(N__4629),
            .I(N__4620));
    LocalMux I__1024 (
            .O(N__4626),
            .I(N__4617));
    Span4Mux_h I__1023 (
            .O(N__4623),
            .I(N__4614));
    InMux I__1022 (
            .O(N__4620),
            .I(N__4611));
    Odrv4 I__1021 (
            .O(N__4617),
            .I(un34_r_val_0_cry_6_c_RNI3LIVZ0));
    Odrv4 I__1020 (
            .O(N__4614),
            .I(un34_r_val_0_cry_6_c_RNI3LIVZ0));
    LocalMux I__1019 (
            .O(N__4611),
            .I(un34_r_val_0_cry_6_c_RNI3LIVZ0));
    InMux I__1018 (
            .O(N__4604),
            .I(N__4594));
    InMux I__1017 (
            .O(N__4603),
            .I(N__4594));
    InMux I__1016 (
            .O(N__4602),
            .I(N__4589));
    InMux I__1015 (
            .O(N__4601),
            .I(N__4589));
    CascadeMux I__1014 (
            .O(N__4600),
            .I(N__4585));
    InMux I__1013 (
            .O(N__4599),
            .I(N__4580));
    LocalMux I__1012 (
            .O(N__4594),
            .I(N__4577));
    LocalMux I__1011 (
            .O(N__4589),
            .I(N__4574));
    InMux I__1010 (
            .O(N__4588),
            .I(N__4569));
    InMux I__1009 (
            .O(N__4585),
            .I(N__4569));
    InMux I__1008 (
            .O(N__4584),
            .I(N__4566));
    InMux I__1007 (
            .O(N__4583),
            .I(N__4563));
    LocalMux I__1006 (
            .O(N__4580),
            .I(N__4560));
    Span4Mux_h I__1005 (
            .O(N__4577),
            .I(N__4557));
    Span4Mux_h I__1004 (
            .O(N__4574),
            .I(N__4552));
    LocalMux I__1003 (
            .O(N__4569),
            .I(N__4552));
    LocalMux I__1002 (
            .O(N__4566),
            .I(ctrZ0Z_25));
    LocalMux I__1001 (
            .O(N__4563),
            .I(ctrZ0Z_25));
    Odrv4 I__1000 (
            .O(N__4560),
            .I(ctrZ0Z_25));
    Odrv4 I__999 (
            .O(N__4557),
            .I(ctrZ0Z_25));
    Odrv4 I__998 (
            .O(N__4552),
            .I(ctrZ0Z_25));
    InMux I__997 (
            .O(N__4541),
            .I(N__4536));
    CascadeMux I__996 (
            .O(N__4540),
            .I(N__4529));
    InMux I__995 (
            .O(N__4539),
            .I(N__4525));
    LocalMux I__994 (
            .O(N__4536),
            .I(N__4522));
    InMux I__993 (
            .O(N__4535),
            .I(N__4517));
    InMux I__992 (
            .O(N__4534),
            .I(N__4517));
    CascadeMux I__991 (
            .O(N__4533),
            .I(N__4514));
    InMux I__990 (
            .O(N__4532),
            .I(N__4509));
    InMux I__989 (
            .O(N__4529),
            .I(N__4509));
    InMux I__988 (
            .O(N__4528),
            .I(N__4505));
    LocalMux I__987 (
            .O(N__4525),
            .I(N__4498));
    Span4Mux_v I__986 (
            .O(N__4522),
            .I(N__4498));
    LocalMux I__985 (
            .O(N__4517),
            .I(N__4498));
    InMux I__984 (
            .O(N__4514),
            .I(N__4495));
    LocalMux I__983 (
            .O(N__4509),
            .I(N__4492));
    InMux I__982 (
            .O(N__4508),
            .I(N__4489));
    LocalMux I__981 (
            .O(N__4505),
            .I(N__4484));
    Span4Mux_s2_v I__980 (
            .O(N__4498),
            .I(N__4484));
    LocalMux I__979 (
            .O(N__4495),
            .I(N__4479));
    Span4Mux_v I__978 (
            .O(N__4492),
            .I(N__4479));
    LocalMux I__977 (
            .O(N__4489),
            .I(ctrZ0Z_27));
    Odrv4 I__976 (
            .O(N__4484),
            .I(ctrZ0Z_27));
    Odrv4 I__975 (
            .O(N__4479),
            .I(ctrZ0Z_27));
    CascadeMux I__974 (
            .O(N__4472),
            .I(N__4466));
    InMux I__973 (
            .O(N__4471),
            .I(N__4453));
    InMux I__972 (
            .O(N__4470),
            .I(N__4453));
    InMux I__971 (
            .O(N__4469),
            .I(N__4448));
    InMux I__970 (
            .O(N__4466),
            .I(N__4448));
    InMux I__969 (
            .O(N__4465),
            .I(N__4443));
    InMux I__968 (
            .O(N__4464),
            .I(N__4443));
    CascadeMux I__967 (
            .O(N__4463),
            .I(N__4436));
    InMux I__966 (
            .O(N__4462),
            .I(N__4427));
    InMux I__965 (
            .O(N__4461),
            .I(N__4427));
    InMux I__964 (
            .O(N__4460),
            .I(N__4427));
    InMux I__963 (
            .O(N__4459),
            .I(N__4420));
    InMux I__962 (
            .O(N__4458),
            .I(N__4415));
    LocalMux I__961 (
            .O(N__4453),
            .I(N__4407));
    LocalMux I__960 (
            .O(N__4448),
            .I(N__4402));
    LocalMux I__959 (
            .O(N__4443),
            .I(N__4402));
    InMux I__958 (
            .O(N__4442),
            .I(N__4391));
    InMux I__957 (
            .O(N__4441),
            .I(N__4391));
    InMux I__956 (
            .O(N__4440),
            .I(N__4391));
    InMux I__955 (
            .O(N__4439),
            .I(N__4391));
    InMux I__954 (
            .O(N__4436),
            .I(N__4391));
    InMux I__953 (
            .O(N__4435),
            .I(N__4386));
    InMux I__952 (
            .O(N__4434),
            .I(N__4386));
    LocalMux I__951 (
            .O(N__4427),
            .I(N__4383));
    InMux I__950 (
            .O(N__4426),
            .I(N__4378));
    InMux I__949 (
            .O(N__4425),
            .I(N__4378));
    InMux I__948 (
            .O(N__4424),
            .I(N__4371));
    InMux I__947 (
            .O(N__4423),
            .I(N__4371));
    LocalMux I__946 (
            .O(N__4420),
            .I(N__4368));
    InMux I__945 (
            .O(N__4419),
            .I(N__4363));
    InMux I__944 (
            .O(N__4418),
            .I(N__4363));
    LocalMux I__943 (
            .O(N__4415),
            .I(N__4358));
    CascadeMux I__942 (
            .O(N__4414),
            .I(N__4354));
    CascadeMux I__941 (
            .O(N__4413),
            .I(N__4350));
    InMux I__940 (
            .O(N__4412),
            .I(N__4341));
    InMux I__939 (
            .O(N__4411),
            .I(N__4341));
    InMux I__938 (
            .O(N__4410),
            .I(N__4341));
    Span4Mux_s3_v I__937 (
            .O(N__4407),
            .I(N__4334));
    Span4Mux_s3_v I__936 (
            .O(N__4402),
            .I(N__4334));
    LocalMux I__935 (
            .O(N__4391),
            .I(N__4334));
    LocalMux I__934 (
            .O(N__4386),
            .I(N__4327));
    Span4Mux_v I__933 (
            .O(N__4383),
            .I(N__4327));
    LocalMux I__932 (
            .O(N__4378),
            .I(N__4327));
    InMux I__931 (
            .O(N__4377),
            .I(N__4324));
    InMux I__930 (
            .O(N__4376),
            .I(N__4321));
    LocalMux I__929 (
            .O(N__4371),
            .I(N__4318));
    Span4Mux_s2_v I__928 (
            .O(N__4368),
            .I(N__4313));
    LocalMux I__927 (
            .O(N__4363),
            .I(N__4313));
    InMux I__926 (
            .O(N__4362),
            .I(N__4308));
    InMux I__925 (
            .O(N__4361),
            .I(N__4308));
    Span4Mux_h I__924 (
            .O(N__4358),
            .I(N__4305));
    InMux I__923 (
            .O(N__4357),
            .I(N__4292));
    InMux I__922 (
            .O(N__4354),
            .I(N__4292));
    InMux I__921 (
            .O(N__4353),
            .I(N__4292));
    InMux I__920 (
            .O(N__4350),
            .I(N__4292));
    InMux I__919 (
            .O(N__4349),
            .I(N__4292));
    InMux I__918 (
            .O(N__4348),
            .I(N__4292));
    LocalMux I__917 (
            .O(N__4341),
            .I(N__4287));
    Span4Mux_h I__916 (
            .O(N__4334),
            .I(N__4287));
    Span4Mux_h I__915 (
            .O(N__4327),
            .I(N__4284));
    LocalMux I__914 (
            .O(N__4324),
            .I(ctrZ0Z_31));
    LocalMux I__913 (
            .O(N__4321),
            .I(ctrZ0Z_31));
    Odrv4 I__912 (
            .O(N__4318),
            .I(ctrZ0Z_31));
    Odrv4 I__911 (
            .O(N__4313),
            .I(ctrZ0Z_31));
    LocalMux I__910 (
            .O(N__4308),
            .I(ctrZ0Z_31));
    Odrv4 I__909 (
            .O(N__4305),
            .I(ctrZ0Z_31));
    LocalMux I__908 (
            .O(N__4292),
            .I(ctrZ0Z_31));
    Odrv4 I__907 (
            .O(N__4287),
            .I(ctrZ0Z_31));
    Odrv4 I__906 (
            .O(N__4284),
            .I(ctrZ0Z_31));
    CascadeMux I__905 (
            .O(N__4265),
            .I(N_70_cascade_));
    CascadeMux I__904 (
            .O(N__4262),
            .I(N__4250));
    CascadeMux I__903 (
            .O(N__4261),
            .I(N__4246));
    CascadeMux I__902 (
            .O(N__4260),
            .I(N__4236));
    CascadeMux I__901 (
            .O(N__4259),
            .I(N__4229));
    CascadeMux I__900 (
            .O(N__4258),
            .I(N__4218));
    InMux I__899 (
            .O(N__4257),
            .I(N__4210));
    InMux I__898 (
            .O(N__4256),
            .I(N__4210));
    InMux I__897 (
            .O(N__4255),
            .I(N__4210));
    CascadeMux I__896 (
            .O(N__4254),
            .I(N__4206));
    InMux I__895 (
            .O(N__4253),
            .I(N__4190));
    InMux I__894 (
            .O(N__4250),
            .I(N__4190));
    InMux I__893 (
            .O(N__4249),
            .I(N__4190));
    InMux I__892 (
            .O(N__4246),
            .I(N__4190));
    InMux I__891 (
            .O(N__4245),
            .I(N__4190));
    InMux I__890 (
            .O(N__4244),
            .I(N__4190));
    InMux I__889 (
            .O(N__4243),
            .I(N__4190));
    InMux I__888 (
            .O(N__4242),
            .I(N__4177));
    InMux I__887 (
            .O(N__4241),
            .I(N__4177));
    InMux I__886 (
            .O(N__4240),
            .I(N__4177));
    InMux I__885 (
            .O(N__4239),
            .I(N__4177));
    InMux I__884 (
            .O(N__4236),
            .I(N__4177));
    InMux I__883 (
            .O(N__4235),
            .I(N__4177));
    InMux I__882 (
            .O(N__4234),
            .I(N__4164));
    InMux I__881 (
            .O(N__4233),
            .I(N__4164));
    InMux I__880 (
            .O(N__4232),
            .I(N__4164));
    InMux I__879 (
            .O(N__4229),
            .I(N__4164));
    InMux I__878 (
            .O(N__4228),
            .I(N__4164));
    InMux I__877 (
            .O(N__4227),
            .I(N__4164));
    CascadeMux I__876 (
            .O(N__4226),
            .I(N__4156));
    CascadeMux I__875 (
            .O(N__4225),
            .I(N__4153));
    CascadeMux I__874 (
            .O(N__4224),
            .I(N__4146));
    InMux I__873 (
            .O(N__4223),
            .I(N__4139));
    InMux I__872 (
            .O(N__4222),
            .I(N__4139));
    InMux I__871 (
            .O(N__4221),
            .I(N__4134));
    InMux I__870 (
            .O(N__4218),
            .I(N__4134));
    InMux I__869 (
            .O(N__4217),
            .I(N__4131));
    LocalMux I__868 (
            .O(N__4210),
            .I(N__4128));
    InMux I__867 (
            .O(N__4209),
            .I(N__4121));
    InMux I__866 (
            .O(N__4206),
            .I(N__4121));
    InMux I__865 (
            .O(N__4205),
            .I(N__4121));
    LocalMux I__864 (
            .O(N__4190),
            .I(N__4114));
    LocalMux I__863 (
            .O(N__4177),
            .I(N__4114));
    LocalMux I__862 (
            .O(N__4164),
            .I(N__4114));
    InMux I__861 (
            .O(N__4163),
            .I(N__4107));
    InMux I__860 (
            .O(N__4162),
            .I(N__4107));
    InMux I__859 (
            .O(N__4161),
            .I(N__4107));
    InMux I__858 (
            .O(N__4160),
            .I(N__4104));
    InMux I__857 (
            .O(N__4159),
            .I(N__4097));
    InMux I__856 (
            .O(N__4156),
            .I(N__4097));
    InMux I__855 (
            .O(N__4153),
            .I(N__4097));
    CascadeMux I__854 (
            .O(N__4152),
            .I(N__4092));
    InMux I__853 (
            .O(N__4151),
            .I(N__4083));
    InMux I__852 (
            .O(N__4150),
            .I(N__4083));
    InMux I__851 (
            .O(N__4149),
            .I(N__4083));
    InMux I__850 (
            .O(N__4146),
            .I(N__4076));
    InMux I__849 (
            .O(N__4145),
            .I(N__4076));
    InMux I__848 (
            .O(N__4144),
            .I(N__4076));
    LocalMux I__847 (
            .O(N__4139),
            .I(N__4073));
    LocalMux I__846 (
            .O(N__4134),
            .I(N__4070));
    LocalMux I__845 (
            .O(N__4131),
            .I(N__4059));
    Span4Mux_v I__844 (
            .O(N__4128),
            .I(N__4050));
    LocalMux I__843 (
            .O(N__4121),
            .I(N__4050));
    Span4Mux_v I__842 (
            .O(N__4114),
            .I(N__4050));
    LocalMux I__841 (
            .O(N__4107),
            .I(N__4050));
    LocalMux I__840 (
            .O(N__4104),
            .I(N__4045));
    LocalMux I__839 (
            .O(N__4097),
            .I(N__4045));
    InMux I__838 (
            .O(N__4096),
            .I(N__4034));
    InMux I__837 (
            .O(N__4095),
            .I(N__4034));
    InMux I__836 (
            .O(N__4092),
            .I(N__4034));
    InMux I__835 (
            .O(N__4091),
            .I(N__4034));
    InMux I__834 (
            .O(N__4090),
            .I(N__4034));
    LocalMux I__833 (
            .O(N__4083),
            .I(N__4025));
    LocalMux I__832 (
            .O(N__4076),
            .I(N__4025));
    Span4Mux_h I__831 (
            .O(N__4073),
            .I(N__4025));
    Span4Mux_h I__830 (
            .O(N__4070),
            .I(N__4025));
    InMux I__829 (
            .O(N__4069),
            .I(N__4008));
    InMux I__828 (
            .O(N__4068),
            .I(N__4008));
    InMux I__827 (
            .O(N__4067),
            .I(N__4008));
    InMux I__826 (
            .O(N__4066),
            .I(N__4008));
    InMux I__825 (
            .O(N__4065),
            .I(N__4008));
    InMux I__824 (
            .O(N__4064),
            .I(N__4008));
    InMux I__823 (
            .O(N__4063),
            .I(N__4008));
    InMux I__822 (
            .O(N__4062),
            .I(N__4008));
    Span4Mux_h I__821 (
            .O(N__4059),
            .I(N__4003));
    Span4Mux_h I__820 (
            .O(N__4050),
            .I(N__4003));
    Odrv4 I__819 (
            .O(N__4045),
            .I(ctrZ0Z_30));
    LocalMux I__818 (
            .O(N__4034),
            .I(ctrZ0Z_30));
    Odrv4 I__817 (
            .O(N__4025),
            .I(ctrZ0Z_30));
    LocalMux I__816 (
            .O(N__4008),
            .I(ctrZ0Z_30));
    Odrv4 I__815 (
            .O(N__4003),
            .I(ctrZ0Z_30));
    InMux I__814 (
            .O(N__3992),
            .I(N__3989));
    LocalMux I__813 (
            .O(N__3989),
            .I(pwm_b_1_7));
    CascadeMux I__812 (
            .O(N__3986),
            .I(N__3982));
    InMux I__811 (
            .O(N__3985),
            .I(N__3978));
    InMux I__810 (
            .O(N__3982),
            .I(N__3975));
    InMux I__809 (
            .O(N__3981),
            .I(N__3968));
    LocalMux I__808 (
            .O(N__3978),
            .I(N__3965));
    LocalMux I__807 (
            .O(N__3975),
            .I(N__3962));
    InMux I__806 (
            .O(N__3974),
            .I(N__3957));
    InMux I__805 (
            .O(N__3973),
            .I(N__3957));
    CascadeMux I__804 (
            .O(N__3972),
            .I(N__3953));
    InMux I__803 (
            .O(N__3971),
            .I(N__3949));
    LocalMux I__802 (
            .O(N__3968),
            .I(N__3946));
    Span4Mux_s2_v I__801 (
            .O(N__3965),
            .I(N__3943));
    Span4Mux_h I__800 (
            .O(N__3962),
            .I(N__3938));
    LocalMux I__799 (
            .O(N__3957),
            .I(N__3938));
    InMux I__798 (
            .O(N__3956),
            .I(N__3931));
    InMux I__797 (
            .O(N__3953),
            .I(N__3931));
    InMux I__796 (
            .O(N__3952),
            .I(N__3931));
    LocalMux I__795 (
            .O(N__3949),
            .I(ctrZ0Z_29));
    Odrv4 I__794 (
            .O(N__3946),
            .I(ctrZ0Z_29));
    Odrv4 I__793 (
            .O(N__3943),
            .I(ctrZ0Z_29));
    Odrv4 I__792 (
            .O(N__3938),
            .I(ctrZ0Z_29));
    LocalMux I__791 (
            .O(N__3931),
            .I(ctrZ0Z_29));
    InMux I__790 (
            .O(N__3920),
            .I(N__3917));
    LocalMux I__789 (
            .O(N__3917),
            .I(pwm_r_1_cry_11_c_RNOZ0Z_0));
    CascadeMux I__788 (
            .O(N__3914),
            .I(N__3911));
    InMux I__787 (
            .O(N__3911),
            .I(N__3908));
    LocalMux I__786 (
            .O(N__3908),
            .I(pwm_r_1_11));
    InMux I__785 (
            .O(N__3905),
            .I(N__3902));
    LocalMux I__784 (
            .O(N__3902),
            .I(N__3899));
    Span4Mux_s3_v I__783 (
            .O(N__3899),
            .I(N__3896));
    Odrv4 I__782 (
            .O(N__3896),
            .I(pwm_g_1_6));
    InMux I__781 (
            .O(N__3893),
            .I(N__3890));
    LocalMux I__780 (
            .O(N__3890),
            .I(N__3886));
    InMux I__779 (
            .O(N__3889),
            .I(N__3883));
    Span4Mux_s3_v I__778 (
            .O(N__3886),
            .I(N__3877));
    LocalMux I__777 (
            .O(N__3883),
            .I(N__3877));
    CascadeMux I__776 (
            .O(N__3882),
            .I(N__3874));
    Span4Mux_h I__775 (
            .O(N__3877),
            .I(N__3871));
    InMux I__774 (
            .O(N__3874),
            .I(N__3868));
    Odrv4 I__773 (
            .O(N__3871),
            .I(un34_r_val_0_cry_7_c_RNI6PJVZ0));
    LocalMux I__772 (
            .O(N__3868),
            .I(un34_r_val_0_cry_7_c_RNI6PJVZ0));
    InMux I__771 (
            .O(N__3863),
            .I(N__3860));
    LocalMux I__770 (
            .O(N__3860),
            .I(un33_r_val_cry_7_THRU_CO));
    CascadeMux I__769 (
            .O(N__3857),
            .I(N_95_cascade_));
    CascadeMux I__768 (
            .O(N__3854),
            .I(N__3851));
    InMux I__767 (
            .O(N__3851),
            .I(N__3848));
    LocalMux I__766 (
            .O(N__3848),
            .I(pwm_r_1_8));
    InMux I__765 (
            .O(N__3845),
            .I(N__3842));
    LocalMux I__764 (
            .O(N__3842),
            .I(N__3837));
    InMux I__763 (
            .O(N__3841),
            .I(N__3834));
    CascadeMux I__762 (
            .O(N__3840),
            .I(N__3831));
    Span4Mux_v I__761 (
            .O(N__3837),
            .I(N__3828));
    LocalMux I__760 (
            .O(N__3834),
            .I(N__3825));
    InMux I__759 (
            .O(N__3831),
            .I(N__3822));
    Odrv4 I__758 (
            .O(N__3828),
            .I(un34_r_val_0_cry_5_c_RNI0HHVZ0));
    Odrv4 I__757 (
            .O(N__3825),
            .I(un34_r_val_0_cry_5_c_RNI0HHVZ0));
    LocalMux I__756 (
            .O(N__3822),
            .I(un34_r_val_0_cry_5_c_RNI0HHVZ0));
    CascadeMux I__755 (
            .O(N__3815),
            .I(N_69_cascade_));
    InMux I__754 (
            .O(N__3812),
            .I(N__3808));
    CascadeMux I__753 (
            .O(N__3811),
            .I(N__3800));
    LocalMux I__752 (
            .O(N__3808),
            .I(N__3797));
    InMux I__751 (
            .O(N__3807),
            .I(N__3790));
    InMux I__750 (
            .O(N__3806),
            .I(N__3790));
    InMux I__749 (
            .O(N__3805),
            .I(N__3790));
    CascadeMux I__748 (
            .O(N__3804),
            .I(N__3786));
    InMux I__747 (
            .O(N__3803),
            .I(N__3782));
    InMux I__746 (
            .O(N__3800),
            .I(N__3779));
    Span4Mux_v I__745 (
            .O(N__3797),
            .I(N__3774));
    LocalMux I__744 (
            .O(N__3790),
            .I(N__3774));
    InMux I__743 (
            .O(N__3789),
            .I(N__3769));
    InMux I__742 (
            .O(N__3786),
            .I(N__3769));
    InMux I__741 (
            .O(N__3785),
            .I(N__3766));
    LocalMux I__740 (
            .O(N__3782),
            .I(N__3763));
    LocalMux I__739 (
            .O(N__3779),
            .I(N__3758));
    Span4Mux_h I__738 (
            .O(N__3774),
            .I(N__3758));
    LocalMux I__737 (
            .O(N__3769),
            .I(N__3755));
    LocalMux I__736 (
            .O(N__3766),
            .I(ctrZ0Z_26));
    Odrv4 I__735 (
            .O(N__3763),
            .I(ctrZ0Z_26));
    Odrv4 I__734 (
            .O(N__3758),
            .I(ctrZ0Z_26));
    Odrv4 I__733 (
            .O(N__3755),
            .I(ctrZ0Z_26));
    InMux I__732 (
            .O(N__3746),
            .I(N__3743));
    LocalMux I__731 (
            .O(N__3743),
            .I(N__3740));
    Odrv4 I__730 (
            .O(N__3740),
            .I(pwm_b_1_6));
    CascadeMux I__729 (
            .O(N__3737),
            .I(N__3732));
    InMux I__728 (
            .O(N__3736),
            .I(N__3725));
    InMux I__727 (
            .O(N__3735),
            .I(N__3725));
    InMux I__726 (
            .O(N__3732),
            .I(N__3719));
    InMux I__725 (
            .O(N__3731),
            .I(N__3713));
    InMux I__724 (
            .O(N__3730),
            .I(N__3713));
    LocalMux I__723 (
            .O(N__3725),
            .I(N__3710));
    InMux I__722 (
            .O(N__3724),
            .I(N__3707));
    CascadeMux I__721 (
            .O(N__3723),
            .I(N__3704));
    InMux I__720 (
            .O(N__3722),
            .I(N__3701));
    LocalMux I__719 (
            .O(N__3719),
            .I(N__3698));
    InMux I__718 (
            .O(N__3718),
            .I(N__3695));
    LocalMux I__717 (
            .O(N__3713),
            .I(N__3692));
    Span4Mux_v I__716 (
            .O(N__3710),
            .I(N__3687));
    LocalMux I__715 (
            .O(N__3707),
            .I(N__3687));
    InMux I__714 (
            .O(N__3704),
            .I(N__3684));
    LocalMux I__713 (
            .O(N__3701),
            .I(N__3679));
    Span4Mux_h I__712 (
            .O(N__3698),
            .I(N__3679));
    LocalMux I__711 (
            .O(N__3695),
            .I(ctrZ0Z_28));
    Odrv4 I__710 (
            .O(N__3692),
            .I(ctrZ0Z_28));
    Odrv4 I__709 (
            .O(N__3687),
            .I(ctrZ0Z_28));
    LocalMux I__708 (
            .O(N__3684),
            .I(ctrZ0Z_28));
    Odrv4 I__707 (
            .O(N__3679),
            .I(ctrZ0Z_28));
    InMux I__706 (
            .O(N__3668),
            .I(N__3665));
    LocalMux I__705 (
            .O(N__3665),
            .I(pwm_r_1_cry_10_c_RNOZ0Z_0));
    InMux I__704 (
            .O(N__3662),
            .I(N__3659));
    LocalMux I__703 (
            .O(N__3659),
            .I(pwm_r_1_10));
    InMux I__702 (
            .O(N__3656),
            .I(N__3653));
    LocalMux I__701 (
            .O(N__3653),
            .I(N__3649));
    CascadeMux I__700 (
            .O(N__3652),
            .I(N__3645));
    Span4Mux_v I__699 (
            .O(N__3649),
            .I(N__3642));
    InMux I__698 (
            .O(N__3648),
            .I(N__3639));
    InMux I__697 (
            .O(N__3645),
            .I(N__3636));
    Odrv4 I__696 (
            .O(N__3642),
            .I(un34_r_val_0_cry_3_c_RNIQ8FVZ0));
    LocalMux I__695 (
            .O(N__3639),
            .I(un34_r_val_0_cry_3_c_RNIQ8FVZ0));
    LocalMux I__694 (
            .O(N__3636),
            .I(un34_r_val_0_cry_3_c_RNIQ8FVZ0));
    CascadeMux I__693 (
            .O(N__3629),
            .I(N_67_cascade_));
    CascadeMux I__692 (
            .O(N__3626),
            .I(N__3623));
    InMux I__691 (
            .O(N__3623),
            .I(N__3620));
    LocalMux I__690 (
            .O(N__3620),
            .I(N__3617));
    Odrv4 I__689 (
            .O(N__3617),
            .I(pwm_r_1_2));
    InMux I__688 (
            .O(N__3614),
            .I(N__3610));
    InMux I__687 (
            .O(N__3613),
            .I(N__3607));
    LocalMux I__686 (
            .O(N__3610),
            .I(N__3600));
    LocalMux I__685 (
            .O(N__3607),
            .I(N__3600));
    CascadeMux I__684 (
            .O(N__3606),
            .I(N__3592));
    InMux I__683 (
            .O(N__3605),
            .I(N__3589));
    Span4Mux_h I__682 (
            .O(N__3600),
            .I(N__3586));
    InMux I__681 (
            .O(N__3599),
            .I(N__3583));
    InMux I__680 (
            .O(N__3598),
            .I(N__3576));
    InMux I__679 (
            .O(N__3597),
            .I(N__3576));
    InMux I__678 (
            .O(N__3596),
            .I(N__3576));
    InMux I__677 (
            .O(N__3595),
            .I(N__3571));
    InMux I__676 (
            .O(N__3592),
            .I(N__3571));
    LocalMux I__675 (
            .O(N__3589),
            .I(ctrZ0Z_21));
    Odrv4 I__674 (
            .O(N__3586),
            .I(ctrZ0Z_21));
    LocalMux I__673 (
            .O(N__3583),
            .I(ctrZ0Z_21));
    LocalMux I__672 (
            .O(N__3576),
            .I(ctrZ0Z_21));
    LocalMux I__671 (
            .O(N__3571),
            .I(ctrZ0Z_21));
    InMux I__670 (
            .O(N__3560),
            .I(N__3557));
    LocalMux I__669 (
            .O(N__3557),
            .I(N__3552));
    CascadeMux I__668 (
            .O(N__3556),
            .I(N__3549));
    InMux I__667 (
            .O(N__3555),
            .I(N__3546));
    Span4Mux_h I__666 (
            .O(N__3552),
            .I(N__3543));
    InMux I__665 (
            .O(N__3549),
            .I(N__3540));
    LocalMux I__664 (
            .O(N__3546),
            .I(un34_r_val_0_cry_2_c_RNIN4EVZ0));
    Odrv4 I__663 (
            .O(N__3543),
            .I(un34_r_val_0_cry_2_c_RNIN4EVZ0));
    LocalMux I__662 (
            .O(N__3540),
            .I(un34_r_val_0_cry_2_c_RNIN4EVZ0));
    InMux I__661 (
            .O(N__3533),
            .I(N__3530));
    LocalMux I__660 (
            .O(N__3530),
            .I(un33_r_val_cry_2_THRU_CO));
    CascadeMux I__659 (
            .O(N__3527),
            .I(N_90_cascade_));
    CascadeMux I__658 (
            .O(N__3524),
            .I(N__3521));
    InMux I__657 (
            .O(N__3521),
            .I(N__3518));
    LocalMux I__656 (
            .O(N__3518),
            .I(N__3515));
    Odrv4 I__655 (
            .O(N__3515),
            .I(pwm_r_1_3));
    InMux I__654 (
            .O(N__3512),
            .I(N__3509));
    LocalMux I__653 (
            .O(N__3509),
            .I(un33_r_val_cry_5_THRU_CO));
    CascadeMux I__652 (
            .O(N__3506),
            .I(N_93_cascade_));
    CascadeMux I__651 (
            .O(N__3503),
            .I(N__3500));
    InMux I__650 (
            .O(N__3500),
            .I(N__3497));
    LocalMux I__649 (
            .O(N__3497),
            .I(pwm_r_1_6));
    InMux I__648 (
            .O(N__3494),
            .I(N__3490));
    CascadeMux I__647 (
            .O(N__3493),
            .I(N__3485));
    LocalMux I__646 (
            .O(N__3490),
            .I(N__3482));
    InMux I__645 (
            .O(N__3489),
            .I(N__3479));
    CascadeMux I__644 (
            .O(N__3488),
            .I(N__3474));
    InMux I__643 (
            .O(N__3485),
            .I(N__3469));
    Span4Mux_v I__642 (
            .O(N__3482),
            .I(N__3464));
    LocalMux I__641 (
            .O(N__3479),
            .I(N__3464));
    CascadeMux I__640 (
            .O(N__3478),
            .I(N__3460));
    InMux I__639 (
            .O(N__3477),
            .I(N__3457));
    InMux I__638 (
            .O(N__3474),
            .I(N__3454));
    InMux I__637 (
            .O(N__3473),
            .I(N__3449));
    InMux I__636 (
            .O(N__3472),
            .I(N__3449));
    LocalMux I__635 (
            .O(N__3469),
            .I(N__3446));
    Span4Mux_h I__634 (
            .O(N__3464),
            .I(N__3443));
    InMux I__633 (
            .O(N__3463),
            .I(N__3438));
    InMux I__632 (
            .O(N__3460),
            .I(N__3438));
    LocalMux I__631 (
            .O(N__3457),
            .I(ctrZ0Z_23));
    LocalMux I__630 (
            .O(N__3454),
            .I(ctrZ0Z_23));
    LocalMux I__629 (
            .O(N__3449),
            .I(ctrZ0Z_23));
    Odrv4 I__628 (
            .O(N__3446),
            .I(ctrZ0Z_23));
    Odrv4 I__627 (
            .O(N__3443),
            .I(ctrZ0Z_23));
    LocalMux I__626 (
            .O(N__3438),
            .I(ctrZ0Z_23));
    InMux I__625 (
            .O(N__3425),
            .I(N__3421));
    CascadeMux I__624 (
            .O(N__3424),
            .I(N__3417));
    LocalMux I__623 (
            .O(N__3421),
            .I(N__3414));
    InMux I__622 (
            .O(N__3420),
            .I(N__3411));
    InMux I__621 (
            .O(N__3417),
            .I(N__3408));
    Odrv4 I__620 (
            .O(N__3414),
            .I(un34_r_val_0_cry_4_c_RNITCGVZ0));
    LocalMux I__619 (
            .O(N__3411),
            .I(un34_r_val_0_cry_4_c_RNITCGVZ0));
    LocalMux I__618 (
            .O(N__3408),
            .I(un34_r_val_0_cry_4_c_RNITCGVZ0));
    CascadeMux I__617 (
            .O(N__3401),
            .I(N_68_cascade_));
    InMux I__616 (
            .O(N__3398),
            .I(N__3395));
    LocalMux I__615 (
            .O(N__3395),
            .I(N__3392));
    Span4Mux_h I__614 (
            .O(N__3392),
            .I(N__3389));
    Odrv4 I__613 (
            .O(N__3389),
            .I(pwm_b_1_5));
    CascadeMux I__612 (
            .O(N__3386),
            .I(N__3383));
    InMux I__611 (
            .O(N__3383),
            .I(N__3380));
    LocalMux I__610 (
            .O(N__3380),
            .I(un33_r_val_cry_6_THRU_CO));
    CascadeMux I__609 (
            .O(N__3377),
            .I(N_94_cascade_));
    CascadeMux I__608 (
            .O(N__3374),
            .I(N__3371));
    InMux I__607 (
            .O(N__3371),
            .I(N__3368));
    LocalMux I__606 (
            .O(N__3368),
            .I(pwm_r_1_7));
    InMux I__605 (
            .O(N__3365),
            .I(N__3362));
    LocalMux I__604 (
            .O(N__3362),
            .I(pwm_b_1_8));
    InMux I__603 (
            .O(N__3359),
            .I(N__3355));
    CascadeMux I__602 (
            .O(N__3358),
            .I(N__3352));
    LocalMux I__601 (
            .O(N__3355),
            .I(N__3348));
    InMux I__600 (
            .O(N__3352),
            .I(N__3345));
    InMux I__599 (
            .O(N__3351),
            .I(N__3342));
    Odrv4 I__598 (
            .O(N__3348),
            .I(pwm_ctr_i_8));
    LocalMux I__597 (
            .O(N__3345),
            .I(pwm_ctr_i_8));
    LocalMux I__596 (
            .O(N__3342),
            .I(pwm_ctr_i_8));
    InMux I__595 (
            .O(N__3335),
            .I(N__3331));
    CascadeMux I__594 (
            .O(N__3334),
            .I(N__3328));
    LocalMux I__593 (
            .O(N__3331),
            .I(N__3324));
    InMux I__592 (
            .O(N__3328),
            .I(N__3321));
    InMux I__591 (
            .O(N__3327),
            .I(N__3318));
    Odrv4 I__590 (
            .O(N__3324),
            .I(pwm_ctr_i_9));
    LocalMux I__589 (
            .O(N__3321),
            .I(pwm_ctr_i_9));
    LocalMux I__588 (
            .O(N__3318),
            .I(pwm_ctr_i_9));
    InMux I__587 (
            .O(N__3311),
            .I(N__3308));
    LocalMux I__586 (
            .O(N__3308),
            .I(N__3305));
    Odrv12 I__585 (
            .O(N__3305),
            .I(pwm_b_1_10));
    CascadeMux I__584 (
            .O(N__3302),
            .I(N__3298));
    CascadeMux I__583 (
            .O(N__3301),
            .I(N__3295));
    InMux I__582 (
            .O(N__3298),
            .I(N__3292));
    InMux I__581 (
            .O(N__3295),
            .I(N__3289));
    LocalMux I__580 (
            .O(N__3292),
            .I(N__3285));
    LocalMux I__579 (
            .O(N__3289),
            .I(N__3282));
    InMux I__578 (
            .O(N__3288),
            .I(N__3279));
    Odrv4 I__577 (
            .O(N__3285),
            .I(pwm_ctr_i_10));
    Odrv4 I__576 (
            .O(N__3282),
            .I(pwm_ctr_i_10));
    LocalMux I__575 (
            .O(N__3279),
            .I(pwm_ctr_i_10));
    InMux I__574 (
            .O(N__3272),
            .I(N__3269));
    LocalMux I__573 (
            .O(N__3269),
            .I(N__3266));
    Odrv4 I__572 (
            .O(N__3266),
            .I(pwm_b_1_11));
    CascadeMux I__571 (
            .O(N__3263),
            .I(N__3259));
    InMux I__570 (
            .O(N__3262),
            .I(N__3256));
    InMux I__569 (
            .O(N__3259),
            .I(N__3253));
    LocalMux I__568 (
            .O(N__3256),
            .I(N__3249));
    LocalMux I__567 (
            .O(N__3253),
            .I(N__3246));
    InMux I__566 (
            .O(N__3252),
            .I(N__3243));
    Odrv4 I__565 (
            .O(N__3249),
            .I(pwm_ctr_i_11));
    Odrv4 I__564 (
            .O(N__3246),
            .I(pwm_ctr_i_11));
    LocalMux I__563 (
            .O(N__3243),
            .I(pwm_ctr_i_11));
    InMux I__562 (
            .O(N__3236),
            .I(pwm_b_1));
    InMux I__561 (
            .O(N__3233),
            .I(N__3230));
    LocalMux I__560 (
            .O(N__3230),
            .I(N__3227));
    Odrv4 I__559 (
            .O(N__3227),
            .I(pwm_bZ0));
    ClkMux I__558 (
            .O(N__3224),
            .I(N__3197));
    ClkMux I__557 (
            .O(N__3223),
            .I(N__3197));
    ClkMux I__556 (
            .O(N__3222),
            .I(N__3197));
    ClkMux I__555 (
            .O(N__3221),
            .I(N__3197));
    ClkMux I__554 (
            .O(N__3220),
            .I(N__3197));
    ClkMux I__553 (
            .O(N__3219),
            .I(N__3197));
    ClkMux I__552 (
            .O(N__3218),
            .I(N__3197));
    ClkMux I__551 (
            .O(N__3217),
            .I(N__3197));
    ClkMux I__550 (
            .O(N__3216),
            .I(N__3197));
    GlobalMux I__549 (
            .O(N__3197),
            .I(clk));
    InMux I__548 (
            .O(N__3194),
            .I(N__3191));
    LocalMux I__547 (
            .O(N__3191),
            .I(N__3187));
    CascadeMux I__546 (
            .O(N__3190),
            .I(N__3183));
    Span4Mux_s1_v I__545 (
            .O(N__3187),
            .I(N__3180));
    InMux I__544 (
            .O(N__3186),
            .I(N__3177));
    InMux I__543 (
            .O(N__3183),
            .I(N__3174));
    Odrv4 I__542 (
            .O(N__3180),
            .I(un34_r_val_0_cry_8_c_RNI9TKVZ0));
    LocalMux I__541 (
            .O(N__3177),
            .I(un34_r_val_0_cry_8_c_RNI9TKVZ0));
    LocalMux I__540 (
            .O(N__3174),
            .I(un34_r_val_0_cry_8_c_RNI9TKVZ0));
    CascadeMux I__539 (
            .O(N__3167),
            .I(N_72_cascade_));
    InMux I__538 (
            .O(N__3164),
            .I(N__3161));
    LocalMux I__537 (
            .O(N__3161),
            .I(pwm_b_1_9));
    InMux I__536 (
            .O(N__3158),
            .I(N__3155));
    LocalMux I__535 (
            .O(N__3155),
            .I(un33_r_val_cry_1_THRU_CO));
    CascadeMux I__534 (
            .O(N__3152),
            .I(N_89_cascade_));
    CascadeMux I__533 (
            .O(N__3149),
            .I(N__3145));
    CascadeMux I__532 (
            .O(N__3148),
            .I(N__3142));
    InMux I__531 (
            .O(N__3145),
            .I(N__3138));
    InMux I__530 (
            .O(N__3142),
            .I(N__3135));
    InMux I__529 (
            .O(N__3141),
            .I(N__3132));
    LocalMux I__528 (
            .O(N__3138),
            .I(N__3129));
    LocalMux I__527 (
            .O(N__3135),
            .I(pwm_ctr_i_0));
    LocalMux I__526 (
            .O(N__3132),
            .I(pwm_ctr_i_0));
    Odrv4 I__525 (
            .O(N__3129),
            .I(pwm_ctr_i_0));
    CascadeMux I__524 (
            .O(N__3122),
            .I(N__3118));
    CascadeMux I__523 (
            .O(N__3121),
            .I(N__3115));
    InMux I__522 (
            .O(N__3118),
            .I(N__3112));
    InMux I__521 (
            .O(N__3115),
            .I(N__3108));
    LocalMux I__520 (
            .O(N__3112),
            .I(N__3105));
    InMux I__519 (
            .O(N__3111),
            .I(N__3102));
    LocalMux I__518 (
            .O(N__3108),
            .I(N__3097));
    Span4Mux_h I__517 (
            .O(N__3105),
            .I(N__3097));
    LocalMux I__516 (
            .O(N__3102),
            .I(pwm_ctr_i_1));
    Odrv4 I__515 (
            .O(N__3097),
            .I(pwm_ctr_i_1));
    CascadeMux I__514 (
            .O(N__3092),
            .I(N__3089));
    InMux I__513 (
            .O(N__3089),
            .I(N__3086));
    LocalMux I__512 (
            .O(N__3086),
            .I(pwm_b_1_1));
    InMux I__511 (
            .O(N__3083),
            .I(N__3079));
    CascadeMux I__510 (
            .O(N__3082),
            .I(N__3076));
    LocalMux I__509 (
            .O(N__3079),
            .I(N__3072));
    InMux I__508 (
            .O(N__3076),
            .I(N__3069));
    InMux I__507 (
            .O(N__3075),
            .I(N__3066));
    Odrv4 I__506 (
            .O(N__3072),
            .I(pwm_ctr_i_2));
    LocalMux I__505 (
            .O(N__3069),
            .I(pwm_ctr_i_2));
    LocalMux I__504 (
            .O(N__3066),
            .I(pwm_ctr_i_2));
    InMux I__503 (
            .O(N__3059),
            .I(N__3056));
    LocalMux I__502 (
            .O(N__3056),
            .I(N__3053));
    Odrv4 I__501 (
            .O(N__3053),
            .I(pwm_b_1_3));
    InMux I__500 (
            .O(N__3050),
            .I(N__3046));
    CascadeMux I__499 (
            .O(N__3049),
            .I(N__3043));
    LocalMux I__498 (
            .O(N__3046),
            .I(N__3039));
    InMux I__497 (
            .O(N__3043),
            .I(N__3036));
    InMux I__496 (
            .O(N__3042),
            .I(N__3033));
    Odrv4 I__495 (
            .O(N__3039),
            .I(pwm_ctr_i_3));
    LocalMux I__494 (
            .O(N__3036),
            .I(pwm_ctr_i_3));
    LocalMux I__493 (
            .O(N__3033),
            .I(pwm_ctr_i_3));
    InMux I__492 (
            .O(N__3026),
            .I(N__3023));
    LocalMux I__491 (
            .O(N__3023),
            .I(N__3019));
    CascadeMux I__490 (
            .O(N__3022),
            .I(N__3016));
    Span4Mux_h I__489 (
            .O(N__3019),
            .I(N__3012));
    InMux I__488 (
            .O(N__3016),
            .I(N__3009));
    InMux I__487 (
            .O(N__3015),
            .I(N__3006));
    Odrv4 I__486 (
            .O(N__3012),
            .I(pwm_ctr_i_4));
    LocalMux I__485 (
            .O(N__3009),
            .I(pwm_ctr_i_4));
    LocalMux I__484 (
            .O(N__3006),
            .I(pwm_ctr_i_4));
    InMux I__483 (
            .O(N__2999),
            .I(N__2995));
    CascadeMux I__482 (
            .O(N__2998),
            .I(N__2992));
    LocalMux I__481 (
            .O(N__2995),
            .I(N__2988));
    InMux I__480 (
            .O(N__2992),
            .I(N__2985));
    InMux I__479 (
            .O(N__2991),
            .I(N__2982));
    Odrv4 I__478 (
            .O(N__2988),
            .I(pwm_ctr_i_5));
    LocalMux I__477 (
            .O(N__2985),
            .I(pwm_ctr_i_5));
    LocalMux I__476 (
            .O(N__2982),
            .I(pwm_ctr_i_5));
    InMux I__475 (
            .O(N__2975),
            .I(N__2970));
    CascadeMux I__474 (
            .O(N__2974),
            .I(N__2967));
    CascadeMux I__473 (
            .O(N__2973),
            .I(N__2964));
    LocalMux I__472 (
            .O(N__2970),
            .I(N__2961));
    InMux I__471 (
            .O(N__2967),
            .I(N__2958));
    InMux I__470 (
            .O(N__2964),
            .I(N__2955));
    Span4Mux_h I__469 (
            .O(N__2961),
            .I(N__2952));
    LocalMux I__468 (
            .O(N__2958),
            .I(pwm_ctr_i_6));
    LocalMux I__467 (
            .O(N__2955),
            .I(pwm_ctr_i_6));
    Odrv4 I__466 (
            .O(N__2952),
            .I(pwm_ctr_i_6));
    InMux I__465 (
            .O(N__2945),
            .I(N__2941));
    CascadeMux I__464 (
            .O(N__2944),
            .I(N__2938));
    LocalMux I__463 (
            .O(N__2941),
            .I(N__2935));
    InMux I__462 (
            .O(N__2938),
            .I(N__2932));
    Span4Mux_h I__461 (
            .O(N__2935),
            .I(N__2928));
    LocalMux I__460 (
            .O(N__2932),
            .I(N__2925));
    InMux I__459 (
            .O(N__2931),
            .I(N__2922));
    Odrv4 I__458 (
            .O(N__2928),
            .I(pwm_ctr_i_7));
    Odrv4 I__457 (
            .O(N__2925),
            .I(pwm_ctr_i_7));
    LocalMux I__456 (
            .O(N__2922),
            .I(pwm_ctr_i_7));
    InMux I__455 (
            .O(N__2915),
            .I(pwm_r_1));
    InMux I__454 (
            .O(N__2912),
            .I(N__2909));
    LocalMux I__453 (
            .O(N__2909),
            .I(N__2906));
    Span4Mux_s2_v I__452 (
            .O(N__2906),
            .I(N__2903));
    Odrv4 I__451 (
            .O(N__2903),
            .I(pwm_rZ0));
    InMux I__450 (
            .O(N__2900),
            .I(N__2897));
    LocalMux I__449 (
            .O(N__2897),
            .I(N__2894));
    Odrv4 I__448 (
            .O(N__2894),
            .I(un33_r_val_cry_8_THRU_CO));
    CascadeMux I__447 (
            .O(N__2891),
            .I(N_96_cascade_));
    CascadeMux I__446 (
            .O(N__2888),
            .I(N__2885));
    InMux I__445 (
            .O(N__2885),
            .I(N__2882));
    LocalMux I__444 (
            .O(N__2882),
            .I(pwm_r_1_9));
    CascadeMux I__443 (
            .O(N__2879),
            .I(N__2875));
    InMux I__442 (
            .O(N__2878),
            .I(N__2872));
    InMux I__441 (
            .O(N__2875),
            .I(N__2869));
    LocalMux I__440 (
            .O(N__2872),
            .I(un34_r_val_0_cry_9_c_RNIV0HKZ0));
    LocalMux I__439 (
            .O(N__2869),
            .I(un34_r_val_0_cry_9_c_RNIV0HKZ0));
    InMux I__438 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__437 (
            .O(N__2861),
            .I(un33_r_val_cry_3_THRU_CO));
    CascadeMux I__436 (
            .O(N__2858),
            .I(N_91_cascade_));
    InMux I__435 (
            .O(N__2855),
            .I(N__2852));
    LocalMux I__434 (
            .O(N__2852),
            .I(pwm_r_1_0));
    InMux I__433 (
            .O(N__2849),
            .I(N__2846));
    LocalMux I__432 (
            .O(N__2846),
            .I(N__2843));
    Odrv4 I__431 (
            .O(N__2843),
            .I(pwm_r_1_1));
    CascadeMux I__430 (
            .O(N__2840),
            .I(N__2837));
    InMux I__429 (
            .O(N__2837),
            .I(N__2834));
    LocalMux I__428 (
            .O(N__2834),
            .I(pwm_r_1_4));
    CascadeMux I__427 (
            .O(N__2831),
            .I(N__2828));
    InMux I__426 (
            .O(N__2828),
            .I(N__2825));
    LocalMux I__425 (
            .O(N__2825),
            .I(pwm_r_1_5));
    InMux I__424 (
            .O(N__2822),
            .I(un33_r_val_cry_3));
    InMux I__423 (
            .O(N__2819),
            .I(N__2816));
    LocalMux I__422 (
            .O(N__2816),
            .I(N__2813));
    Odrv4 I__421 (
            .O(N__2813),
            .I(un33_r_val_cry_4_THRU_CO));
    InMux I__420 (
            .O(N__2810),
            .I(un33_r_val_cry_4));
    InMux I__419 (
            .O(N__2807),
            .I(un33_r_val_cry_5));
    InMux I__418 (
            .O(N__2804),
            .I(un33_r_val_cry_6));
    InMux I__417 (
            .O(N__2801),
            .I(bfn_3_26_0_));
    InMux I__416 (
            .O(N__2798),
            .I(N__2795));
    LocalMux I__415 (
            .O(N__2795),
            .I(N__2791));
    InMux I__414 (
            .O(N__2794),
            .I(N__2787));
    Span4Mux_v I__413 (
            .O(N__2791),
            .I(N__2783));
    InMux I__412 (
            .O(N__2790),
            .I(N__2780));
    LocalMux I__411 (
            .O(N__2787),
            .I(N__2777));
    InMux I__410 (
            .O(N__2786),
            .I(N__2774));
    Sp12to4 I__409 (
            .O(N__2783),
            .I(N__2770));
    LocalMux I__408 (
            .O(N__2780),
            .I(N__2763));
    Span4Mux_s1_v I__407 (
            .O(N__2777),
            .I(N__2763));
    LocalMux I__406 (
            .O(N__2774),
            .I(N__2763));
    CascadeMux I__405 (
            .O(N__2773),
            .I(N__2752));
    Span12Mux_h I__404 (
            .O(N__2770),
            .I(N__2749));
    Span4Mux_v I__403 (
            .O(N__2763),
            .I(N__2746));
    InMux I__402 (
            .O(N__2762),
            .I(N__2743));
    InMux I__401 (
            .O(N__2761),
            .I(N__2740));
    InMux I__400 (
            .O(N__2760),
            .I(N__2733));
    InMux I__399 (
            .O(N__2759),
            .I(N__2733));
    InMux I__398 (
            .O(N__2758),
            .I(N__2733));
    InMux I__397 (
            .O(N__2757),
            .I(N__2724));
    InMux I__396 (
            .O(N__2756),
            .I(N__2724));
    InMux I__395 (
            .O(N__2755),
            .I(N__2724));
    InMux I__394 (
            .O(N__2752),
            .I(N__2724));
    Odrv12 I__393 (
            .O(N__2749),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__392 (
            .O(N__2746),
            .I(CONSTANT_ONE_NET));
    LocalMux I__391 (
            .O(N__2743),
            .I(CONSTANT_ONE_NET));
    LocalMux I__390 (
            .O(N__2740),
            .I(CONSTANT_ONE_NET));
    LocalMux I__389 (
            .O(N__2733),
            .I(CONSTANT_ONE_NET));
    LocalMux I__388 (
            .O(N__2724),
            .I(CONSTANT_ONE_NET));
    InMux I__387 (
            .O(N__2711),
            .I(un33_r_val_cry_8));
    InMux I__386 (
            .O(N__2708),
            .I(un33_r_val_cry_9));
    InMux I__385 (
            .O(N__2705),
            .I(un33_r_val_cry_10));
    CascadeMux I__384 (
            .O(N__2702),
            .I(un33_r_val_cry_10_THRU_CO_cascade_));
    InMux I__383 (
            .O(N__2699),
            .I(N__2696));
    LocalMux I__382 (
            .O(N__2696),
            .I(un34_r_val_0_cry_10_THRU_CO));
    CascadeMux I__381 (
            .O(N__2693),
            .I(N__2690));
    InMux I__380 (
            .O(N__2690),
            .I(N__2687));
    LocalMux I__379 (
            .O(N__2687),
            .I(N__2684));
    Odrv4 I__378 (
            .O(N__2684),
            .I(pwm_g_1_11));
    InMux I__377 (
            .O(N__2681),
            .I(pwm_g_1));
    InMux I__376 (
            .O(N__2678),
            .I(N__2675));
    LocalMux I__375 (
            .O(N__2675),
            .I(N__2672));
    Odrv4 I__374 (
            .O(N__2672),
            .I(pwm_gZ0));
    CascadeMux I__373 (
            .O(N__2669),
            .I(N_71_cascade_));
    CascadeMux I__372 (
            .O(N__2666),
            .I(N__2663));
    InMux I__371 (
            .O(N__2663),
            .I(N__2660));
    LocalMux I__370 (
            .O(N__2660),
            .I(pwm_g_1_10));
    InMux I__369 (
            .O(N__2657),
            .I(N__2653));
    InMux I__368 (
            .O(N__2656),
            .I(N__2650));
    LocalMux I__367 (
            .O(N__2653),
            .I(ctr_RNI7D9MZ0Z_21));
    LocalMux I__366 (
            .O(N__2650),
            .I(ctr_RNI7D9MZ0Z_21));
    InMux I__365 (
            .O(N__2645),
            .I(N__2642));
    LocalMux I__364 (
            .O(N__2642),
            .I(un33_r_val_cry_0_THRU_CO));
    InMux I__363 (
            .O(N__2639),
            .I(un33_r_val_cry_0));
    InMux I__362 (
            .O(N__2636),
            .I(un33_r_val_cry_1));
    InMux I__361 (
            .O(N__2633),
            .I(un33_r_val_cry_2));
    InMux I__360 (
            .O(N__2630),
            .I(N__2626));
    InMux I__359 (
            .O(N__2629),
            .I(N__2623));
    LocalMux I__358 (
            .O(N__2626),
            .I(pwm_ctrZ0Z_3));
    LocalMux I__357 (
            .O(N__2623),
            .I(pwm_ctrZ0Z_3));
    CascadeMux I__356 (
            .O(N__2618),
            .I(N__2615));
    InMux I__355 (
            .O(N__2615),
            .I(N__2612));
    LocalMux I__354 (
            .O(N__2612),
            .I(pwm_g_1_3));
    InMux I__353 (
            .O(N__2609),
            .I(N__2605));
    InMux I__352 (
            .O(N__2608),
            .I(N__2602));
    LocalMux I__351 (
            .O(N__2605),
            .I(pwm_ctrZ0Z_4));
    LocalMux I__350 (
            .O(N__2602),
            .I(pwm_ctrZ0Z_4));
    CascadeMux I__349 (
            .O(N__2597),
            .I(N__2594));
    InMux I__348 (
            .O(N__2594),
            .I(N__2591));
    LocalMux I__347 (
            .O(N__2591),
            .I(N__2588));
    Span4Mux_s2_v I__346 (
            .O(N__2588),
            .I(N__2585));
    Odrv4 I__345 (
            .O(N__2585),
            .I(pwm_g_1_5));
    InMux I__344 (
            .O(N__2582),
            .I(N__2578));
    InMux I__343 (
            .O(N__2581),
            .I(N__2575));
    LocalMux I__342 (
            .O(N__2578),
            .I(pwm_ctrZ0Z_5));
    LocalMux I__341 (
            .O(N__2575),
            .I(pwm_ctrZ0Z_5));
    InMux I__340 (
            .O(N__2570),
            .I(N__2566));
    InMux I__339 (
            .O(N__2569),
            .I(N__2563));
    LocalMux I__338 (
            .O(N__2566),
            .I(pwm_ctrZ0Z_6));
    LocalMux I__337 (
            .O(N__2563),
            .I(pwm_ctrZ0Z_6));
    InMux I__336 (
            .O(N__2558),
            .I(N__2554));
    InMux I__335 (
            .O(N__2557),
            .I(N__2551));
    LocalMux I__334 (
            .O(N__2554),
            .I(pwm_ctrZ0Z_7));
    LocalMux I__333 (
            .O(N__2551),
            .I(pwm_ctrZ0Z_7));
    CascadeMux I__332 (
            .O(N__2546),
            .I(N__2543));
    InMux I__331 (
            .O(N__2543),
            .I(N__2540));
    LocalMux I__330 (
            .O(N__2540),
            .I(pwm_g_1_8));
    InMux I__329 (
            .O(N__2537),
            .I(N__2533));
    InMux I__328 (
            .O(N__2536),
            .I(N__2530));
    LocalMux I__327 (
            .O(N__2533),
            .I(pwm_ctrZ0Z_8));
    LocalMux I__326 (
            .O(N__2530),
            .I(pwm_ctrZ0Z_8));
    CascadeMux I__325 (
            .O(N__2525),
            .I(N__2522));
    InMux I__324 (
            .O(N__2522),
            .I(N__2519));
    LocalMux I__323 (
            .O(N__2519),
            .I(N__2516));
    Odrv4 I__322 (
            .O(N__2516),
            .I(pwm_g_1_9));
    InMux I__321 (
            .O(N__2513),
            .I(N__2509));
    InMux I__320 (
            .O(N__2512),
            .I(N__2506));
    LocalMux I__319 (
            .O(N__2509),
            .I(pwm_ctrZ0Z_9));
    LocalMux I__318 (
            .O(N__2506),
            .I(pwm_ctrZ0Z_9));
    InMux I__317 (
            .O(N__2501),
            .I(N__2497));
    InMux I__316 (
            .O(N__2500),
            .I(N__2494));
    LocalMux I__315 (
            .O(N__2497),
            .I(pwm_ctrZ0Z_10));
    LocalMux I__314 (
            .O(N__2494),
            .I(pwm_ctrZ0Z_10));
    InMux I__313 (
            .O(N__2489),
            .I(N__2485));
    InMux I__312 (
            .O(N__2488),
            .I(N__2482));
    LocalMux I__311 (
            .O(N__2485),
            .I(pwm_ctrZ0Z_11));
    LocalMux I__310 (
            .O(N__2482),
            .I(pwm_ctrZ0Z_11));
    CascadeMux I__309 (
            .O(N__2477),
            .I(N_87_cascade_));
    CascadeMux I__308 (
            .O(N__2474),
            .I(N__2471));
    InMux I__307 (
            .O(N__2471),
            .I(N__2468));
    LocalMux I__306 (
            .O(N__2468),
            .I(N__2462));
    InMux I__305 (
            .O(N__2467),
            .I(N__2459));
    InMux I__304 (
            .O(N__2466),
            .I(N__2454));
    InMux I__303 (
            .O(N__2465),
            .I(N__2454));
    Span4Mux_v I__302 (
            .O(N__2462),
            .I(N__2451));
    LocalMux I__301 (
            .O(N__2459),
            .I(ctrZ0Z_19));
    LocalMux I__300 (
            .O(N__2454),
            .I(ctrZ0Z_19));
    Odrv4 I__299 (
            .O(N__2451),
            .I(ctrZ0Z_19));
    CascadeMux I__298 (
            .O(N__2444),
            .I(un40_b_val_3_ns_1_1_cascade_));
    CascadeMux I__297 (
            .O(N__2441),
            .I(N__2438));
    InMux I__296 (
            .O(N__2438),
            .I(N__2435));
    LocalMux I__295 (
            .O(N__2435),
            .I(pwm_g_1_0));
    InMux I__294 (
            .O(N__2432),
            .I(N__2428));
    InMux I__293 (
            .O(N__2431),
            .I(N__2425));
    LocalMux I__292 (
            .O(N__2428),
            .I(pwm_ctrZ0Z_0));
    LocalMux I__291 (
            .O(N__2425),
            .I(pwm_ctrZ0Z_0));
    InMux I__290 (
            .O(N__2420),
            .I(N__2416));
    InMux I__289 (
            .O(N__2419),
            .I(N__2413));
    LocalMux I__288 (
            .O(N__2416),
            .I(pwm_ctrZ0Z_1));
    LocalMux I__287 (
            .O(N__2413),
            .I(pwm_ctrZ0Z_1));
    InMux I__286 (
            .O(N__2408),
            .I(N__2405));
    LocalMux I__285 (
            .O(N__2405),
            .I(pwm_g_1_1));
    InMux I__284 (
            .O(N__2402),
            .I(N__2398));
    InMux I__283 (
            .O(N__2401),
            .I(N__2395));
    LocalMux I__282 (
            .O(N__2398),
            .I(pwm_ctrZ0Z_2));
    LocalMux I__281 (
            .O(N__2395),
            .I(pwm_ctrZ0Z_2));
    CascadeMux I__280 (
            .O(N__2390),
            .I(N__2387));
    InMux I__279 (
            .O(N__2387),
            .I(N__2384));
    LocalMux I__278 (
            .O(N__2384),
            .I(pwm_g_1_2));
    InMux I__277 (
            .O(N__2381),
            .I(un34_r_val_0_cry_9));
    InMux I__276 (
            .O(N__2378),
            .I(un34_r_val_0_cry_10));
    CascadeMux I__275 (
            .O(N__2375),
            .I(un34_r_val_0_cry_10_THRU_CO_cascade_));
    CascadeMux I__274 (
            .O(N__2372),
            .I(N_92_cascade_));
    CascadeMux I__273 (
            .O(N__2369),
            .I(N_66_cascade_));
    InMux I__272 (
            .O(N__2366),
            .I(un34_r_val_0_cry_1));
    InMux I__271 (
            .O(N__2363),
            .I(un34_r_val_0_cry_2));
    InMux I__270 (
            .O(N__2360),
            .I(un34_r_val_0_cry_3));
    InMux I__269 (
            .O(N__2357),
            .I(un34_r_val_0_cry_4));
    InMux I__268 (
            .O(N__2354),
            .I(un34_r_val_0_cry_5));
    InMux I__267 (
            .O(N__2351),
            .I(un34_r_val_0_cry_6));
    InMux I__266 (
            .O(N__2348),
            .I(un34_r_val_0_cry_7));
    InMux I__265 (
            .O(N__2345),
            .I(bfn_2_27_0_));
    InMux I__264 (
            .O(N__2342),
            .I(pwm_ctr_cry_8));
    InMux I__263 (
            .O(N__2339),
            .I(pwm_ctr_cry_9));
    InMux I__262 (
            .O(N__2336),
            .I(pwm_ctr_cry_10));
    CascadeMux I__261 (
            .O(N__2333),
            .I(N_88_cascade_));
    InMux I__260 (
            .O(N__2330),
            .I(bfn_1_29_0_));
    InMux I__259 (
            .O(N__2327),
            .I(pwm_ctr_cry_0));
    InMux I__258 (
            .O(N__2324),
            .I(pwm_ctr_cry_1));
    InMux I__257 (
            .O(N__2321),
            .I(pwm_ctr_cry_2));
    InMux I__256 (
            .O(N__2318),
            .I(pwm_ctr_cry_3));
    InMux I__255 (
            .O(N__2315),
            .I(pwm_ctr_cry_4));
    InMux I__254 (
            .O(N__2312),
            .I(pwm_ctr_cry_5));
    InMux I__253 (
            .O(N__2309),
            .I(pwm_ctr_cry_6));
    InMux I__252 (
            .O(N__2306),
            .I(bfn_1_30_0_));
    InMux I__251 (
            .O(N__2303),
            .I(ctr_cry_22));
    InMux I__250 (
            .O(N__2300),
            .I(bfn_1_28_0_));
    InMux I__249 (
            .O(N__2297),
            .I(ctr_cry_24));
    InMux I__248 (
            .O(N__2294),
            .I(ctr_cry_25));
    InMux I__247 (
            .O(N__2291),
            .I(ctr_cry_26));
    InMux I__246 (
            .O(N__2288),
            .I(ctr_cry_27));
    InMux I__245 (
            .O(N__2285),
            .I(ctr_cry_28));
    InMux I__244 (
            .O(N__2282),
            .I(ctr_cry_29));
    InMux I__243 (
            .O(N__2279),
            .I(ctr_cry_30));
    InMux I__242 (
            .O(N__2276),
            .I(N__2273));
    LocalMux I__241 (
            .O(N__2273),
            .I(ctrZ0Z_14));
    InMux I__240 (
            .O(N__2270),
            .I(ctr_cry_13));
    InMux I__239 (
            .O(N__2267),
            .I(N__2264));
    LocalMux I__238 (
            .O(N__2264),
            .I(ctrZ0Z_15));
    InMux I__237 (
            .O(N__2261),
            .I(ctr_cry_14));
    InMux I__236 (
            .O(N__2258),
            .I(N__2255));
    LocalMux I__235 (
            .O(N__2255),
            .I(ctrZ0Z_16));
    InMux I__234 (
            .O(N__2252),
            .I(bfn_1_27_0_));
    InMux I__233 (
            .O(N__2249),
            .I(N__2246));
    LocalMux I__232 (
            .O(N__2246),
            .I(ctrZ0Z_17));
    InMux I__231 (
            .O(N__2243),
            .I(ctr_cry_16));
    InMux I__230 (
            .O(N__2240),
            .I(ctr_cry_17));
    InMux I__229 (
            .O(N__2237),
            .I(ctr_cry_18));
    InMux I__228 (
            .O(N__2234),
            .I(ctr_cry_19));
    InMux I__227 (
            .O(N__2231),
            .I(ctr_cry_20));
    InMux I__226 (
            .O(N__2228),
            .I(ctr_cry_21));
    InMux I__225 (
            .O(N__2225),
            .I(N__2222));
    LocalMux I__224 (
            .O(N__2222),
            .I(ctrZ0Z_6));
    InMux I__223 (
            .O(N__2219),
            .I(ctr_cry_5));
    InMux I__222 (
            .O(N__2216),
            .I(N__2213));
    LocalMux I__221 (
            .O(N__2213),
            .I(ctrZ0Z_7));
    InMux I__220 (
            .O(N__2210),
            .I(ctr_cry_6));
    InMux I__219 (
            .O(N__2207),
            .I(N__2204));
    LocalMux I__218 (
            .O(N__2204),
            .I(ctrZ0Z_8));
    InMux I__217 (
            .O(N__2201),
            .I(bfn_1_26_0_));
    InMux I__216 (
            .O(N__2198),
            .I(N__2195));
    LocalMux I__215 (
            .O(N__2195),
            .I(ctrZ0Z_9));
    InMux I__214 (
            .O(N__2192),
            .I(ctr_cry_8));
    InMux I__213 (
            .O(N__2189),
            .I(N__2186));
    LocalMux I__212 (
            .O(N__2186),
            .I(ctrZ0Z_10));
    InMux I__211 (
            .O(N__2183),
            .I(ctr_cry_9));
    InMux I__210 (
            .O(N__2180),
            .I(N__2177));
    LocalMux I__209 (
            .O(N__2177),
            .I(ctrZ0Z_11));
    InMux I__208 (
            .O(N__2174),
            .I(ctr_cry_10));
    InMux I__207 (
            .O(N__2171),
            .I(N__2168));
    LocalMux I__206 (
            .O(N__2168),
            .I(ctrZ0Z_12));
    InMux I__205 (
            .O(N__2165),
            .I(ctr_cry_11));
    InMux I__204 (
            .O(N__2162),
            .I(N__2159));
    LocalMux I__203 (
            .O(N__2159),
            .I(ctrZ0Z_13));
    InMux I__202 (
            .O(N__2156),
            .I(ctr_cry_12));
    InMux I__201 (
            .O(N__2153),
            .I(N__2150));
    LocalMux I__200 (
            .O(N__2150),
            .I(ctrZ0Z_0));
    InMux I__199 (
            .O(N__2147),
            .I(bfn_1_25_0_));
    InMux I__198 (
            .O(N__2144),
            .I(N__2141));
    LocalMux I__197 (
            .O(N__2141),
            .I(ctrZ0Z_1));
    InMux I__196 (
            .O(N__2138),
            .I(ctr_cry_0));
    InMux I__195 (
            .O(N__2135),
            .I(N__2132));
    LocalMux I__194 (
            .O(N__2132),
            .I(ctrZ0Z_2));
    InMux I__193 (
            .O(N__2129),
            .I(ctr_cry_1));
    InMux I__192 (
            .O(N__2126),
            .I(N__2123));
    LocalMux I__191 (
            .O(N__2123),
            .I(ctrZ0Z_3));
    InMux I__190 (
            .O(N__2120),
            .I(ctr_cry_2));
    InMux I__189 (
            .O(N__2117),
            .I(N__2114));
    LocalMux I__188 (
            .O(N__2114),
            .I(ctrZ0Z_4));
    InMux I__187 (
            .O(N__2111),
            .I(ctr_cry_3));
    InMux I__186 (
            .O(N__2108),
            .I(N__2105));
    LocalMux I__185 (
            .O(N__2105),
            .I(ctrZ0Z_5));
    InMux I__184 (
            .O(N__2102),
            .I(ctr_cry_4));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(un33_r_val_cry_7),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_3_27_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_27_0_));
    defparam IN_MUX_bfv_3_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_28_0_ (
            .carryinitin(pwm_r_1_cry_7),
            .carryinitout(bfn_3_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_3_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_30_0_ (
            .carryinitin(pwm_b_1_cry_7),
            .carryinitout(bfn_3_30_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(pwm_g_1_cry_7),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_1_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_29_0_));
    defparam IN_MUX_bfv_1_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_30_0_ (
            .carryinitin(pwm_ctr_cry_7),
            .carryinitout(bfn_1_30_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_1_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_26_0_ (
            .carryinitin(ctr_cry_7),
            .carryinitout(bfn_1_26_0_));
    defparam IN_MUX_bfv_1_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_27_0_ (
            .carryinitin(ctr_cry_15),
            .carryinitout(bfn_1_27_0_));
    defparam IN_MUX_bfv_1_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_28_0_ (
            .carryinitin(ctr_cry_23),
            .carryinitout(bfn_1_28_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(un34_r_val_0_cry_8),
            .carryinitout(bfn_2_27_0_));
    VCC VCC (
            .Y(VCCG0));
    defparam RGBA_DRIVER.CURRENT_MODE="0b1";
    defparam RGBA_DRIVER.RGB2_CURRENT="0b000111";
    defparam RGBA_DRIVER.RGB1_CURRENT="0b000111";
    defparam RGBA_DRIVER.RGB0_CURRENT="0b000111";
    SB_RGBA_DRV RGBA_DRIVER (
            .RGBLEDEN(N__2794),
            .RGB2PWM(N__2912),
            .RGB1(RGB1),
            .CURREN(N__2798),
            .RGB2(RGB2),
            .RGB1PWM(N__3233),
            .RGB0PWM(N__2678),
            .RGB0(RGB0));
    defparam inthosc.CLKHF_DIV="0b00";
    SB_HFOSC inthosc (
            .CLKHFPU(N__2786),
            .CLKHFEN(N__2790),
            .CLKHF(clk));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam ctr_0_LC_1_25_0.C_ON=1'b1;
    defparam ctr_0_LC_1_25_0.SEQ_MODE=4'b1000;
    defparam ctr_0_LC_1_25_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_0_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__2153),
            .in2(_gnd_net_),
            .in3(N__2147),
            .lcout(ctrZ0Z_0),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(ctr_cry_0),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_1_LC_1_25_1.C_ON=1'b1;
    defparam ctr_1_LC_1_25_1.SEQ_MODE=4'b1000;
    defparam ctr_1_LC_1_25_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_1_LC_1_25_1 (
            .in0(_gnd_net_),
            .in1(N__2144),
            .in2(_gnd_net_),
            .in3(N__2138),
            .lcout(ctrZ0Z_1),
            .ltout(),
            .carryin(ctr_cry_0),
            .carryout(ctr_cry_1),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_2_LC_1_25_2.C_ON=1'b1;
    defparam ctr_2_LC_1_25_2.SEQ_MODE=4'b1000;
    defparam ctr_2_LC_1_25_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_2_LC_1_25_2 (
            .in0(_gnd_net_),
            .in1(N__2135),
            .in2(_gnd_net_),
            .in3(N__2129),
            .lcout(ctrZ0Z_2),
            .ltout(),
            .carryin(ctr_cry_1),
            .carryout(ctr_cry_2),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_3_LC_1_25_3.C_ON=1'b1;
    defparam ctr_3_LC_1_25_3.SEQ_MODE=4'b1000;
    defparam ctr_3_LC_1_25_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_3_LC_1_25_3 (
            .in0(_gnd_net_),
            .in1(N__2126),
            .in2(_gnd_net_),
            .in3(N__2120),
            .lcout(ctrZ0Z_3),
            .ltout(),
            .carryin(ctr_cry_2),
            .carryout(ctr_cry_3),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_4_LC_1_25_4.C_ON=1'b1;
    defparam ctr_4_LC_1_25_4.SEQ_MODE=4'b1000;
    defparam ctr_4_LC_1_25_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_4_LC_1_25_4 (
            .in0(_gnd_net_),
            .in1(N__2117),
            .in2(_gnd_net_),
            .in3(N__2111),
            .lcout(ctrZ0Z_4),
            .ltout(),
            .carryin(ctr_cry_3),
            .carryout(ctr_cry_4),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_5_LC_1_25_5.C_ON=1'b1;
    defparam ctr_5_LC_1_25_5.SEQ_MODE=4'b1000;
    defparam ctr_5_LC_1_25_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_5_LC_1_25_5 (
            .in0(_gnd_net_),
            .in1(N__2108),
            .in2(_gnd_net_),
            .in3(N__2102),
            .lcout(ctrZ0Z_5),
            .ltout(),
            .carryin(ctr_cry_4),
            .carryout(ctr_cry_5),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_6_LC_1_25_6.C_ON=1'b1;
    defparam ctr_6_LC_1_25_6.SEQ_MODE=4'b1000;
    defparam ctr_6_LC_1_25_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_6_LC_1_25_6 (
            .in0(_gnd_net_),
            .in1(N__2225),
            .in2(_gnd_net_),
            .in3(N__2219),
            .lcout(ctrZ0Z_6),
            .ltout(),
            .carryin(ctr_cry_5),
            .carryout(ctr_cry_6),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_7_LC_1_25_7.C_ON=1'b1;
    defparam ctr_7_LC_1_25_7.SEQ_MODE=4'b1000;
    defparam ctr_7_LC_1_25_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_7_LC_1_25_7 (
            .in0(_gnd_net_),
            .in1(N__2216),
            .in2(_gnd_net_),
            .in3(N__2210),
            .lcout(ctrZ0Z_7),
            .ltout(),
            .carryin(ctr_cry_6),
            .carryout(ctr_cry_7),
            .clk(N__3224),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_8_LC_1_26_0.C_ON=1'b1;
    defparam ctr_8_LC_1_26_0.SEQ_MODE=4'b1000;
    defparam ctr_8_LC_1_26_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_8_LC_1_26_0 (
            .in0(_gnd_net_),
            .in1(N__2207),
            .in2(_gnd_net_),
            .in3(N__2201),
            .lcout(ctrZ0Z_8),
            .ltout(),
            .carryin(bfn_1_26_0_),
            .carryout(ctr_cry_8),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_9_LC_1_26_1.C_ON=1'b1;
    defparam ctr_9_LC_1_26_1.SEQ_MODE=4'b1000;
    defparam ctr_9_LC_1_26_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_9_LC_1_26_1 (
            .in0(_gnd_net_),
            .in1(N__2198),
            .in2(_gnd_net_),
            .in3(N__2192),
            .lcout(ctrZ0Z_9),
            .ltout(),
            .carryin(ctr_cry_8),
            .carryout(ctr_cry_9),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_10_LC_1_26_2.C_ON=1'b1;
    defparam ctr_10_LC_1_26_2.SEQ_MODE=4'b1000;
    defparam ctr_10_LC_1_26_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_10_LC_1_26_2 (
            .in0(_gnd_net_),
            .in1(N__2189),
            .in2(_gnd_net_),
            .in3(N__2183),
            .lcout(ctrZ0Z_10),
            .ltout(),
            .carryin(ctr_cry_9),
            .carryout(ctr_cry_10),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_11_LC_1_26_3.C_ON=1'b1;
    defparam ctr_11_LC_1_26_3.SEQ_MODE=4'b1000;
    defparam ctr_11_LC_1_26_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_11_LC_1_26_3 (
            .in0(_gnd_net_),
            .in1(N__2180),
            .in2(_gnd_net_),
            .in3(N__2174),
            .lcout(ctrZ0Z_11),
            .ltout(),
            .carryin(ctr_cry_10),
            .carryout(ctr_cry_11),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_12_LC_1_26_4.C_ON=1'b1;
    defparam ctr_12_LC_1_26_4.SEQ_MODE=4'b1000;
    defparam ctr_12_LC_1_26_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_12_LC_1_26_4 (
            .in0(_gnd_net_),
            .in1(N__2171),
            .in2(_gnd_net_),
            .in3(N__2165),
            .lcout(ctrZ0Z_12),
            .ltout(),
            .carryin(ctr_cry_11),
            .carryout(ctr_cry_12),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_13_LC_1_26_5.C_ON=1'b1;
    defparam ctr_13_LC_1_26_5.SEQ_MODE=4'b1000;
    defparam ctr_13_LC_1_26_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_13_LC_1_26_5 (
            .in0(_gnd_net_),
            .in1(N__2162),
            .in2(_gnd_net_),
            .in3(N__2156),
            .lcout(ctrZ0Z_13),
            .ltout(),
            .carryin(ctr_cry_12),
            .carryout(ctr_cry_13),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_14_LC_1_26_6.C_ON=1'b1;
    defparam ctr_14_LC_1_26_6.SEQ_MODE=4'b1000;
    defparam ctr_14_LC_1_26_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_14_LC_1_26_6 (
            .in0(_gnd_net_),
            .in1(N__2276),
            .in2(_gnd_net_),
            .in3(N__2270),
            .lcout(ctrZ0Z_14),
            .ltout(),
            .carryin(ctr_cry_13),
            .carryout(ctr_cry_14),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_15_LC_1_26_7.C_ON=1'b1;
    defparam ctr_15_LC_1_26_7.SEQ_MODE=4'b1000;
    defparam ctr_15_LC_1_26_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_15_LC_1_26_7 (
            .in0(_gnd_net_),
            .in1(N__2267),
            .in2(_gnd_net_),
            .in3(N__2261),
            .lcout(ctrZ0Z_15),
            .ltout(),
            .carryin(ctr_cry_14),
            .carryout(ctr_cry_15),
            .clk(N__3222),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_16_LC_1_27_0.C_ON=1'b1;
    defparam ctr_16_LC_1_27_0.SEQ_MODE=4'b1000;
    defparam ctr_16_LC_1_27_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_16_LC_1_27_0 (
            .in0(_gnd_net_),
            .in1(N__2258),
            .in2(_gnd_net_),
            .in3(N__2252),
            .lcout(ctrZ0Z_16),
            .ltout(),
            .carryin(bfn_1_27_0_),
            .carryout(ctr_cry_16),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_17_LC_1_27_1.C_ON=1'b1;
    defparam ctr_17_LC_1_27_1.SEQ_MODE=4'b1000;
    defparam ctr_17_LC_1_27_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_17_LC_1_27_1 (
            .in0(_gnd_net_),
            .in1(N__2249),
            .in2(_gnd_net_),
            .in3(N__2243),
            .lcout(ctrZ0Z_17),
            .ltout(),
            .carryin(ctr_cry_16),
            .carryout(ctr_cry_17),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_18_LC_1_27_2.C_ON=1'b1;
    defparam ctr_18_LC_1_27_2.SEQ_MODE=4'b1000;
    defparam ctr_18_LC_1_27_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_18_LC_1_27_2 (
            .in0(_gnd_net_),
            .in1(N__4938),
            .in2(_gnd_net_),
            .in3(N__2240),
            .lcout(ctrZ0Z_18),
            .ltout(),
            .carryin(ctr_cry_17),
            .carryout(ctr_cry_18),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_19_LC_1_27_3.C_ON=1'b1;
    defparam ctr_19_LC_1_27_3.SEQ_MODE=4'b1000;
    defparam ctr_19_LC_1_27_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_19_LC_1_27_3 (
            .in0(_gnd_net_),
            .in1(N__2467),
            .in2(_gnd_net_),
            .in3(N__2237),
            .lcout(ctrZ0Z_19),
            .ltout(),
            .carryin(ctr_cry_18),
            .carryout(ctr_cry_19),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_20_LC_1_27_4.C_ON=1'b1;
    defparam ctr_20_LC_1_27_4.SEQ_MODE=4'b1000;
    defparam ctr_20_LC_1_27_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_20_LC_1_27_4 (
            .in0(_gnd_net_),
            .in1(N__4852),
            .in2(_gnd_net_),
            .in3(N__2234),
            .lcout(ctrZ0Z_20),
            .ltout(),
            .carryin(ctr_cry_19),
            .carryout(ctr_cry_20),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_21_LC_1_27_5.C_ON=1'b1;
    defparam ctr_21_LC_1_27_5.SEQ_MODE=4'b1000;
    defparam ctr_21_LC_1_27_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_21_LC_1_27_5 (
            .in0(_gnd_net_),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__2231),
            .lcout(ctrZ0Z_21),
            .ltout(),
            .carryin(ctr_cry_20),
            .carryout(ctr_cry_21),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_22_LC_1_27_6.C_ON=1'b1;
    defparam ctr_22_LC_1_27_6.SEQ_MODE=4'b1000;
    defparam ctr_22_LC_1_27_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_22_LC_1_27_6 (
            .in0(_gnd_net_),
            .in1(N__4770),
            .in2(_gnd_net_),
            .in3(N__2228),
            .lcout(ctrZ0Z_22),
            .ltout(),
            .carryin(ctr_cry_21),
            .carryout(ctr_cry_22),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_23_LC_1_27_7.C_ON=1'b1;
    defparam ctr_23_LC_1_27_7.SEQ_MODE=4'b1000;
    defparam ctr_23_LC_1_27_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_23_LC_1_27_7 (
            .in0(_gnd_net_),
            .in1(N__3477),
            .in2(_gnd_net_),
            .in3(N__2303),
            .lcout(ctrZ0Z_23),
            .ltout(),
            .carryin(ctr_cry_22),
            .carryout(ctr_cry_23),
            .clk(N__3221),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_24_LC_1_28_0.C_ON=1'b1;
    defparam ctr_24_LC_1_28_0.SEQ_MODE=4'b1000;
    defparam ctr_24_LC_1_28_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_24_LC_1_28_0 (
            .in0(_gnd_net_),
            .in1(N__4720),
            .in2(_gnd_net_),
            .in3(N__2300),
            .lcout(ctrZ0Z_24),
            .ltout(),
            .carryin(bfn_1_28_0_),
            .carryout(ctr_cry_24),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_25_LC_1_28_1.C_ON=1'b1;
    defparam ctr_25_LC_1_28_1.SEQ_MODE=4'b1000;
    defparam ctr_25_LC_1_28_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_25_LC_1_28_1 (
            .in0(_gnd_net_),
            .in1(N__4584),
            .in2(_gnd_net_),
            .in3(N__2297),
            .lcout(ctrZ0Z_25),
            .ltout(),
            .carryin(ctr_cry_24),
            .carryout(ctr_cry_25),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_26_LC_1_28_2.C_ON=1'b1;
    defparam ctr_26_LC_1_28_2.SEQ_MODE=4'b1000;
    defparam ctr_26_LC_1_28_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_26_LC_1_28_2 (
            .in0(_gnd_net_),
            .in1(N__3785),
            .in2(_gnd_net_),
            .in3(N__2294),
            .lcout(ctrZ0Z_26),
            .ltout(),
            .carryin(ctr_cry_25),
            .carryout(ctr_cry_26),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_27_LC_1_28_3.C_ON=1'b1;
    defparam ctr_27_LC_1_28_3.SEQ_MODE=4'b1000;
    defparam ctr_27_LC_1_28_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_27_LC_1_28_3 (
            .in0(_gnd_net_),
            .in1(N__4508),
            .in2(_gnd_net_),
            .in3(N__2291),
            .lcout(ctrZ0Z_27),
            .ltout(),
            .carryin(ctr_cry_26),
            .carryout(ctr_cry_27),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_28_LC_1_28_4.C_ON=1'b1;
    defparam ctr_28_LC_1_28_4.SEQ_MODE=4'b1000;
    defparam ctr_28_LC_1_28_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_28_LC_1_28_4 (
            .in0(_gnd_net_),
            .in1(N__3718),
            .in2(_gnd_net_),
            .in3(N__2288),
            .lcout(ctrZ0Z_28),
            .ltout(),
            .carryin(ctr_cry_27),
            .carryout(ctr_cry_28),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_29_LC_1_28_5.C_ON=1'b1;
    defparam ctr_29_LC_1_28_5.SEQ_MODE=4'b1000;
    defparam ctr_29_LC_1_28_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_29_LC_1_28_5 (
            .in0(_gnd_net_),
            .in1(N__3971),
            .in2(_gnd_net_),
            .in3(N__2285),
            .lcout(ctrZ0Z_29),
            .ltout(),
            .carryin(ctr_cry_28),
            .carryout(ctr_cry_29),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_30_LC_1_28_6.C_ON=1'b1;
    defparam ctr_30_LC_1_28_6.SEQ_MODE=4'b1000;
    defparam ctr_30_LC_1_28_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 ctr_30_LC_1_28_6 (
            .in0(_gnd_net_),
            .in1(N__4160),
            .in2(_gnd_net_),
            .in3(N__2282),
            .lcout(ctrZ0Z_30),
            .ltout(),
            .carryin(ctr_cry_29),
            .carryout(ctr_cry_30),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_31_LC_1_28_7.C_ON=1'b0;
    defparam ctr_31_LC_1_28_7.SEQ_MODE=4'b1000;
    defparam ctr_31_LC_1_28_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 ctr_31_LC_1_28_7 (
            .in0(_gnd_net_),
            .in1(N__4377),
            .in2(_gnd_net_),
            .in3(N__2279),
            .lcout(ctrZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3219),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_0_LC_1_29_0.C_ON=1'b1;
    defparam pwm_ctr_0_LC_1_29_0.SEQ_MODE=4'b1000;
    defparam pwm_ctr_0_LC_1_29_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_0_LC_1_29_0 (
            .in0(_gnd_net_),
            .in1(N__2432),
            .in2(_gnd_net_),
            .in3(N__2330),
            .lcout(pwm_ctrZ0Z_0),
            .ltout(),
            .carryin(bfn_1_29_0_),
            .carryout(pwm_ctr_cry_0),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_1_LC_1_29_1.C_ON=1'b1;
    defparam pwm_ctr_1_LC_1_29_1.SEQ_MODE=4'b1000;
    defparam pwm_ctr_1_LC_1_29_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_1_LC_1_29_1 (
            .in0(_gnd_net_),
            .in1(N__2420),
            .in2(_gnd_net_),
            .in3(N__2327),
            .lcout(pwm_ctrZ0Z_1),
            .ltout(),
            .carryin(pwm_ctr_cry_0),
            .carryout(pwm_ctr_cry_1),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_2_LC_1_29_2.C_ON=1'b1;
    defparam pwm_ctr_2_LC_1_29_2.SEQ_MODE=4'b1000;
    defparam pwm_ctr_2_LC_1_29_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_2_LC_1_29_2 (
            .in0(_gnd_net_),
            .in1(N__2402),
            .in2(_gnd_net_),
            .in3(N__2324),
            .lcout(pwm_ctrZ0Z_2),
            .ltout(),
            .carryin(pwm_ctr_cry_1),
            .carryout(pwm_ctr_cry_2),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_3_LC_1_29_3.C_ON=1'b1;
    defparam pwm_ctr_3_LC_1_29_3.SEQ_MODE=4'b1000;
    defparam pwm_ctr_3_LC_1_29_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_3_LC_1_29_3 (
            .in0(_gnd_net_),
            .in1(N__2630),
            .in2(_gnd_net_),
            .in3(N__2321),
            .lcout(pwm_ctrZ0Z_3),
            .ltout(),
            .carryin(pwm_ctr_cry_2),
            .carryout(pwm_ctr_cry_3),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_4_LC_1_29_4.C_ON=1'b1;
    defparam pwm_ctr_4_LC_1_29_4.SEQ_MODE=4'b1000;
    defparam pwm_ctr_4_LC_1_29_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_4_LC_1_29_4 (
            .in0(_gnd_net_),
            .in1(N__2609),
            .in2(_gnd_net_),
            .in3(N__2318),
            .lcout(pwm_ctrZ0Z_4),
            .ltout(),
            .carryin(pwm_ctr_cry_3),
            .carryout(pwm_ctr_cry_4),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_5_LC_1_29_5.C_ON=1'b1;
    defparam pwm_ctr_5_LC_1_29_5.SEQ_MODE=4'b1000;
    defparam pwm_ctr_5_LC_1_29_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_5_LC_1_29_5 (
            .in0(_gnd_net_),
            .in1(N__2582),
            .in2(_gnd_net_),
            .in3(N__2315),
            .lcout(pwm_ctrZ0Z_5),
            .ltout(),
            .carryin(pwm_ctr_cry_4),
            .carryout(pwm_ctr_cry_5),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_6_LC_1_29_6.C_ON=1'b1;
    defparam pwm_ctr_6_LC_1_29_6.SEQ_MODE=4'b1000;
    defparam pwm_ctr_6_LC_1_29_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_6_LC_1_29_6 (
            .in0(_gnd_net_),
            .in1(N__2570),
            .in2(_gnd_net_),
            .in3(N__2312),
            .lcout(pwm_ctrZ0Z_6),
            .ltout(),
            .carryin(pwm_ctr_cry_5),
            .carryout(pwm_ctr_cry_6),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_7_LC_1_29_7.C_ON=1'b1;
    defparam pwm_ctr_7_LC_1_29_7.SEQ_MODE=4'b1000;
    defparam pwm_ctr_7_LC_1_29_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_7_LC_1_29_7 (
            .in0(_gnd_net_),
            .in1(N__2558),
            .in2(_gnd_net_),
            .in3(N__2309),
            .lcout(pwm_ctrZ0Z_7),
            .ltout(),
            .carryin(pwm_ctr_cry_6),
            .carryout(pwm_ctr_cry_7),
            .clk(N__3217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_8_LC_1_30_0.C_ON=1'b1;
    defparam pwm_ctr_8_LC_1_30_0.SEQ_MODE=4'b1000;
    defparam pwm_ctr_8_LC_1_30_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_8_LC_1_30_0 (
            .in0(_gnd_net_),
            .in1(N__2537),
            .in2(_gnd_net_),
            .in3(N__2306),
            .lcout(pwm_ctrZ0Z_8),
            .ltout(),
            .carryin(bfn_1_30_0_),
            .carryout(pwm_ctr_cry_8),
            .clk(N__3216),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_9_LC_1_30_1.C_ON=1'b1;
    defparam pwm_ctr_9_LC_1_30_1.SEQ_MODE=4'b1000;
    defparam pwm_ctr_9_LC_1_30_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_9_LC_1_30_1 (
            .in0(_gnd_net_),
            .in1(N__2513),
            .in2(_gnd_net_),
            .in3(N__2342),
            .lcout(pwm_ctrZ0Z_9),
            .ltout(),
            .carryin(pwm_ctr_cry_8),
            .carryout(pwm_ctr_cry_9),
            .clk(N__3216),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_10_LC_1_30_2.C_ON=1'b1;
    defparam pwm_ctr_10_LC_1_30_2.SEQ_MODE=4'b1000;
    defparam pwm_ctr_10_LC_1_30_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 pwm_ctr_10_LC_1_30_2 (
            .in0(_gnd_net_),
            .in1(N__2501),
            .in2(_gnd_net_),
            .in3(N__2339),
            .lcout(pwm_ctrZ0Z_10),
            .ltout(),
            .carryin(pwm_ctr_cry_9),
            .carryout(pwm_ctr_cry_10),
            .clk(N__3216),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctr_11_LC_1_30_3.C_ON=1'b0;
    defparam pwm_ctr_11_LC_1_30_3.SEQ_MODE=4'b1000;
    defparam pwm_ctr_11_LC_1_30_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 pwm_ctr_11_LC_1_30_3 (
            .in0(_gnd_net_),
            .in1(N__2489),
            .in2(_gnd_net_),
            .in3(N__2336),
            .lcout(pwm_ctrZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3216),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIVDLC1_27_LC_1_30_5.C_ON=1'b0;
    defparam ctr_RNIVDLC1_27_LC_1_30_5.SEQ_MODE=4'b0000;
    defparam ctr_RNIVDLC1_27_LC_1_30_5.LUT_INIT=16'b1101100000011011;
    LogicCell40 ctr_RNIVDLC1_27_LC_1_30_5 (
            .in0(N__4410),
            .in1(N__3973),
            .in2(N__4533),
            .in3(N__4150),
            .lcout(pwm_g_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNITBLC1_26_LC_1_30_6.C_ON=1'b0;
    defparam ctr_RNITBLC1_26_LC_1_30_6.SEQ_MODE=4'b0000;
    defparam ctr_RNITBLC1_26_LC_1_30_6.LUT_INIT=16'b1000110110110001;
    LogicCell40 ctr_RNITBLC1_26_LC_1_30_6 (
            .in0(N__4149),
            .in1(N__3722),
            .in2(N__3811),
            .in3(N__4412),
            .lcout(pwm_g_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNILGG11_29_LC_1_30_7.C_ON=1'b0;
    defparam ctr_RNILGG11_29_LC_1_30_7.SEQ_MODE=4'b0000;
    defparam ctr_RNILGG11_29_LC_1_30_7.LUT_INIT=16'b0100010000100010;
    LogicCell40 ctr_RNILGG11_29_LC_1_30_7 (
            .in0(N__4411),
            .in1(N__4151),
            .in2(_gnd_net_),
            .in3(N__3974),
            .lcout(pwm_g_1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_1_c_RNO_0_LC_2_25_1.C_ON=1'b0;
    defparam pwm_r_1_cry_1_c_RNO_0_LC_2_25_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_1_c_RNO_0_LC_2_25_1.LUT_INIT=16'b0100111000011011;
    LogicCell40 pwm_r_1_cry_1_c_RNO_0_LC_2_25_1 (
            .in0(N__4161),
            .in1(N__2657),
            .in2(N__2474),
            .in3(N__2645),
            .lcout(),
            .ltout(N_88_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_1_c_RNO_LC_2_25_2.C_ON=1'b0;
    defparam pwm_r_1_cry_1_c_RNO_LC_2_25_2.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_1_c_RNO_LC_2_25_2.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_1_c_RNO_LC_2_25_2 (
            .in0(N__4425),
            .in1(N__4162),
            .in2(N__2333),
            .in3(N__3614),
            .lcout(pwm_r_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIN5LC1_23_LC_2_25_4.C_ON=1'b0;
    defparam ctr_RNIN5LC1_23_LC_2_25_4.SEQ_MODE=4'b0000;
    defparam ctr_RNIN5LC1_23_LC_2_25_4.LUT_INIT=16'b1101100000011011;
    LogicCell40 ctr_RNIN5LC1_23_LC_2_25_4 (
            .in0(N__4426),
            .in1(N__4599),
            .in2(N__3493),
            .in3(N__4163),
            .lcout(pwm_g_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_25_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_25_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_25_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNI7D9M_21_LC_2_26_0.C_ON=1'b1;
    defparam ctr_RNI7D9M_21_LC_2_26_0.SEQ_MODE=4'b0000;
    defparam ctr_RNI7D9M_21_LC_2_26_0.LUT_INIT=16'b0011110000111100;
    LogicCell40 ctr_RNI7D9M_21_LC_2_26_0 (
            .in0(_gnd_net_),
            .in1(N__4836),
            .in2(N__3606),
            .in3(_gnd_net_),
            .lcout(ctr_RNI7D9MZ0Z_21),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(un34_r_val_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_1_c_RNIK0DV_LC_2_26_1.C_ON=1'b1;
    defparam un34_r_val_0_cry_1_c_RNIK0DV_LC_2_26_1.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_1_c_RNIK0DV_LC_2_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_1_c_RNIK0DV_LC_2_26_1 (
            .in0(_gnd_net_),
            .in1(N__3595),
            .in2(N__4771),
            .in3(N__2366),
            .lcout(un34_r_val_0_cry_1_c_RNIK0DVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_1),
            .carryout(un34_r_val_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_2_c_RNIN4EV_LC_2_26_2.C_ON=1'b1;
    defparam un34_r_val_0_cry_2_c_RNIN4EV_LC_2_26_2.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_2_c_RNIN4EV_LC_2_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_2_c_RNIN4EV_LC_2_26_2 (
            .in0(_gnd_net_),
            .in1(N__4758),
            .in2(N__3478),
            .in3(N__2363),
            .lcout(un34_r_val_0_cry_2_c_RNIN4EVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_2),
            .carryout(un34_r_val_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_3_c_RNIQ8FV_LC_2_26_3.C_ON=1'b1;
    defparam un34_r_val_0_cry_3_c_RNIQ8FV_LC_2_26_3.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_3_c_RNIQ8FV_LC_2_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_3_c_RNIQ8FV_LC_2_26_3 (
            .in0(_gnd_net_),
            .in1(N__3463),
            .in2(N__4721),
            .in3(N__2360),
            .lcout(un34_r_val_0_cry_3_c_RNIQ8FVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_3),
            .carryout(un34_r_val_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_4_c_RNITCGV_LC_2_26_4.C_ON=1'b1;
    defparam un34_r_val_0_cry_4_c_RNITCGV_LC_2_26_4.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_4_c_RNITCGV_LC_2_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_4_c_RNITCGV_LC_2_26_4 (
            .in0(_gnd_net_),
            .in1(N__4702),
            .in2(N__4600),
            .in3(N__2357),
            .lcout(un34_r_val_0_cry_4_c_RNITCGVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_4),
            .carryout(un34_r_val_0_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_5_c_RNI0HHV_LC_2_26_5.C_ON=1'b1;
    defparam un34_r_val_0_cry_5_c_RNI0HHV_LC_2_26_5.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_5_c_RNI0HHV_LC_2_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_5_c_RNI0HHV_LC_2_26_5 (
            .in0(_gnd_net_),
            .in1(N__4588),
            .in2(N__3804),
            .in3(N__2354),
            .lcout(un34_r_val_0_cry_5_c_RNI0HHVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_5),
            .carryout(un34_r_val_0_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_6_c_RNI3LIV_LC_2_26_6.C_ON=1'b1;
    defparam un34_r_val_0_cry_6_c_RNI3LIV_LC_2_26_6.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_6_c_RNI3LIV_LC_2_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_6_c_RNI3LIV_LC_2_26_6 (
            .in0(_gnd_net_),
            .in1(N__3789),
            .in2(N__4540),
            .in3(N__2351),
            .lcout(un34_r_val_0_cry_6_c_RNI3LIVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_6),
            .carryout(un34_r_val_0_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_7_c_RNI6PJV_LC_2_26_7.C_ON=1'b1;
    defparam un34_r_val_0_cry_7_c_RNI6PJV_LC_2_26_7.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_7_c_RNI6PJV_LC_2_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_7_c_RNI6PJV_LC_2_26_7 (
            .in0(_gnd_net_),
            .in1(N__4532),
            .in2(N__3737),
            .in3(N__2348),
            .lcout(un34_r_val_0_cry_7_c_RNI6PJVZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_7),
            .carryout(un34_r_val_0_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_8_c_RNI9TKV_LC_2_27_0.C_ON=1'b1;
    defparam un34_r_val_0_cry_8_c_RNI9TKV_LC_2_27_0.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_8_c_RNI9TKV_LC_2_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un34_r_val_0_cry_8_c_RNI9TKV_LC_2_27_0 (
            .in0(_gnd_net_),
            .in1(N__3952),
            .in2(N__3723),
            .in3(N__2345),
            .lcout(un34_r_val_0_cry_8_c_RNI9TKVZ0),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(un34_r_val_0_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_9_c_RNIV0HK_LC_2_27_1.C_ON=1'b1;
    defparam un34_r_val_0_cry_9_c_RNIV0HK_LC_2_27_1.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_9_c_RNIV0HK_LC_2_27_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un34_r_val_0_cry_9_c_RNIV0HK_LC_2_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3972),
            .in3(N__2381),
            .lcout(un34_r_val_0_cry_9_c_RNIV0HKZ0),
            .ltout(),
            .carryin(un34_r_val_0_cry_9),
            .carryout(un34_r_val_0_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un34_r_val_0_cry_10_THRU_LUT4_0_LC_2_27_2.C_ON=1'b0;
    defparam un34_r_val_0_cry_10_THRU_LUT4_0_LC_2_27_2.SEQ_MODE=4'b0000;
    defparam un34_r_val_0_cry_10_THRU_LUT4_0_LC_2_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un34_r_val_0_cry_10_THRU_LUT4_0_LC_2_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2378),
            .lcout(un34_r_val_0_cry_10_THRU_CO),
            .ltout(un34_r_val_0_cry_10_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_11_c_RNO_LC_2_27_3.C_ON=1'b0;
    defparam pwm_b_1_cry_11_c_RNO_LC_2_27_3.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_11_c_RNO_LC_2_27_3.LUT_INIT=16'b0000110010001000;
    LogicCell40 pwm_b_1_cry_11_c_RNO_LC_2_27_3 (
            .in0(N__3956),
            .in1(N__4376),
            .in2(N__2375),
            .in3(N__4096),
            .lcout(pwm_b_1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_5_c_RNO_0_LC_2_27_4.C_ON=1'b0;
    defparam pwm_r_1_cry_5_c_RNO_0_LC_2_27_4.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_5_c_RNO_0_LC_2_27_4.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_5_c_RNO_0_LC_2_27_4 (
            .in0(N__3472),
            .in1(N__3420),
            .in2(N__4152),
            .in3(N__2819),
            .lcout(),
            .ltout(N_92_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_5_c_RNO_LC_2_27_5.C_ON=1'b0;
    defparam pwm_r_1_cry_5_c_RNO_LC_2_27_5.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_5_c_RNO_LC_2_27_5.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_5_c_RNO_LC_2_27_5 (
            .in0(N__4362),
            .in1(N__4095),
            .in2(N__2372),
            .in3(N__4583),
            .lcout(pwm_r_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_3_c_RNO_0_LC_2_27_6.C_ON=1'b0;
    defparam pwm_b_1_cry_3_c_RNO_0_LC_2_27_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_3_c_RNO_0_LC_2_27_6.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_3_c_RNO_0_LC_2_27_6 (
            .in0(N__4090),
            .in1(N__3599),
            .in2(_gnd_net_),
            .in3(N__3555),
            .lcout(),
            .ltout(N_66_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_3_c_RNO_LC_2_27_7.C_ON=1'b0;
    defparam pwm_b_1_cry_3_c_RNO_LC_2_27_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_3_c_RNO_LC_2_27_7.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_3_c_RNO_LC_2_27_7 (
            .in0(N__4361),
            .in1(N__4091),
            .in2(N__2369),
            .in3(N__3473),
            .lcout(pwm_b_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIO5KC1_19_LC_2_28_0.C_ON=1'b0;
    defparam ctr_RNIO5KC1_19_LC_2_28_0.SEQ_MODE=4'b0000;
    defparam ctr_RNIO5KC1_19_LC_2_28_0.LUT_INIT=16'b1011100000011101;
    LogicCell40 ctr_RNIO5KC1_19_LC_2_28_0 (
            .in0(N__4064),
            .in1(N__2465),
            .in2(N__4413),
            .in3(N__3597),
            .lcout(pwm_g_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIM3KC1_18_LC_2_28_1.C_ON=1'b0;
    defparam ctr_RNIM3KC1_18_LC_2_28_1.SEQ_MODE=4'b0000;
    defparam ctr_RNIM3KC1_18_LC_2_28_1.LUT_INIT=16'b1011100000011101;
    LogicCell40 ctr_RNIM3KC1_18_LC_2_28_1 (
            .in0(N__4850),
            .in1(N__4349),
            .in2(N__4939),
            .in3(N__4066),
            .lcout(pwm_g_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_0_c_RNO_0_LC_2_28_2.C_ON=1'b0;
    defparam pwm_r_1_cry_0_c_RNO_0_LC_2_28_2.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_0_c_RNO_0_LC_2_28_2.LUT_INIT=16'b0010001001110111;
    LogicCell40 pwm_r_1_cry_0_c_RNO_0_LC_2_28_2 (
            .in0(N__4062),
            .in1(N__4931),
            .in2(_gnd_net_),
            .in3(N__4847),
            .lcout(),
            .ltout(N_87_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_0_c_RNO_LC_2_28_3.C_ON=1'b0;
    defparam pwm_r_1_cry_0_c_RNO_LC_2_28_3.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_0_c_RNO_LC_2_28_3.LUT_INIT=16'b1011100000110000;
    LogicCell40 pwm_r_1_cry_0_c_RNO_LC_2_28_3 (
            .in0(N__4849),
            .in1(N__4348),
            .in2(N__2477),
            .in3(N__4065),
            .lcout(pwm_r_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIHVKC1_22_LC_2_28_4.C_ON=1'b0;
    defparam ctr_RNIHVKC1_22_LC_2_28_4.SEQ_MODE=4'b0000;
    defparam ctr_RNIHVKC1_22_LC_2_28_4.LUT_INIT=16'b1000101111010001;
    LogicCell40 ctr_RNIHVKC1_22_LC_2_28_4 (
            .in0(N__4067),
            .in1(N__4769),
            .in2(N__4414),
            .in3(N__4851),
            .lcout(pwm_g_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIJ1LC1_21_LC_2_28_5.C_ON=1'b0;
    defparam ctr_RNIJ1LC1_21_LC_2_28_5.SEQ_MODE=4'b0000;
    defparam ctr_RNIJ1LC1_21_LC_2_28_5.LUT_INIT=16'b1101000110001011;
    LogicCell40 ctr_RNIJ1LC1_21_LC_2_28_5 (
            .in0(N__3598),
            .in1(N__4069),
            .in2(N__3488),
            .in3(N__4357),
            .lcout(pwm_g_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_1_c_RNO_0_LC_2_28_6.C_ON=1'b0;
    defparam pwm_b_1_cry_1_c_RNO_0_LC_2_28_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_1_c_RNO_0_LC_2_28_6.LUT_INIT=16'b0011001110011001;
    LogicCell40 pwm_b_1_cry_1_c_RNO_0_LC_2_28_6 (
            .in0(N__4063),
            .in1(N__3596),
            .in2(_gnd_net_),
            .in3(N__4848),
            .lcout(),
            .ltout(un40_b_val_3_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_1_c_RNO_LC_2_28_7.C_ON=1'b0;
    defparam pwm_b_1_cry_1_c_RNO_LC_2_28_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_1_c_RNO_LC_2_28_7.LUT_INIT=16'b0000110010111000;
    LogicCell40 pwm_b_1_cry_1_c_RNO_LC_2_28_7 (
            .in0(N__2466),
            .in1(N__4353),
            .in2(N__2444),
            .in3(N__4068),
            .lcout(pwm_b_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_0_c_inv_LC_2_29_0.C_ON=1'b1;
    defparam pwm_g_1_cry_0_c_inv_LC_2_29_0.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_0_c_inv_LC_2_29_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_0_c_inv_LC_2_29_0 (
            .in0(_gnd_net_),
            .in1(N__3141),
            .in2(N__2441),
            .in3(N__2431),
            .lcout(pwm_ctr_i_0),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(pwm_g_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_1_c_inv_LC_2_29_1.C_ON=1'b1;
    defparam pwm_g_1_cry_1_c_inv_LC_2_29_1.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_1_c_inv_LC_2_29_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 pwm_g_1_cry_1_c_inv_LC_2_29_1 (
            .in0(N__2419),
            .in1(N__2408),
            .in2(N__3121),
            .in3(_gnd_net_),
            .lcout(pwm_ctr_i_1),
            .ltout(),
            .carryin(pwm_g_1_cry_0),
            .carryout(pwm_g_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_2_c_inv_LC_2_29_2.C_ON=1'b1;
    defparam pwm_g_1_cry_2_c_inv_LC_2_29_2.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_2_c_inv_LC_2_29_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 pwm_g_1_cry_2_c_inv_LC_2_29_2 (
            .in0(N__2401),
            .in1(N__3075),
            .in2(N__2390),
            .in3(_gnd_net_),
            .lcout(pwm_ctr_i_2),
            .ltout(),
            .carryin(pwm_g_1_cry_1),
            .carryout(pwm_g_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_3_c_inv_LC_2_29_3.C_ON=1'b1;
    defparam pwm_g_1_cry_3_c_inv_LC_2_29_3.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_3_c_inv_LC_2_29_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 pwm_g_1_cry_3_c_inv_LC_2_29_3 (
            .in0(N__2629),
            .in1(N__3042),
            .in2(N__2618),
            .in3(_gnd_net_),
            .lcout(pwm_ctr_i_3),
            .ltout(),
            .carryin(pwm_g_1_cry_2),
            .carryout(pwm_g_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_4_c_inv_LC_2_29_4.C_ON=1'b1;
    defparam pwm_g_1_cry_4_c_inv_LC_2_29_4.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_4_c_inv_LC_2_29_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_4_c_inv_LC_2_29_4 (
            .in0(_gnd_net_),
            .in1(N__3015),
            .in2(N__4664),
            .in3(N__2608),
            .lcout(pwm_ctr_i_4),
            .ltout(),
            .carryin(pwm_g_1_cry_3),
            .carryout(pwm_g_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_5_c_inv_LC_2_29_5.C_ON=1'b1;
    defparam pwm_g_1_cry_5_c_inv_LC_2_29_5.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_5_c_inv_LC_2_29_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_5_c_inv_LC_2_29_5 (
            .in0(_gnd_net_),
            .in1(N__2991),
            .in2(N__2597),
            .in3(N__2581),
            .lcout(pwm_ctr_i_5),
            .ltout(),
            .carryin(pwm_g_1_cry_4),
            .carryout(pwm_g_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_6_c_inv_LC_2_29_6.C_ON=1'b1;
    defparam pwm_g_1_cry_6_c_inv_LC_2_29_6.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_6_c_inv_LC_2_29_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_6_c_inv_LC_2_29_6 (
            .in0(_gnd_net_),
            .in1(N__3905),
            .in2(N__2973),
            .in3(N__2569),
            .lcout(pwm_ctr_i_6),
            .ltout(),
            .carryin(pwm_g_1_cry_5),
            .carryout(pwm_g_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_7_c_inv_LC_2_29_7.C_ON=1'b1;
    defparam pwm_g_1_cry_7_c_inv_LC_2_29_7.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_7_c_inv_LC_2_29_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_7_c_inv_LC_2_29_7 (
            .in0(_gnd_net_),
            .in1(N__2931),
            .in2(N__4649),
            .in3(N__2557),
            .lcout(pwm_ctr_i_7),
            .ltout(),
            .carryin(pwm_g_1_cry_6),
            .carryout(pwm_g_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_8_c_inv_LC_2_30_0.C_ON=1'b1;
    defparam pwm_g_1_cry_8_c_inv_LC_2_30_0.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_8_c_inv_LC_2_30_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_8_c_inv_LC_2_30_0 (
            .in0(_gnd_net_),
            .in1(N__3351),
            .in2(N__2546),
            .in3(N__2536),
            .lcout(pwm_ctr_i_8),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(pwm_g_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_9_c_inv_LC_2_30_1.C_ON=1'b1;
    defparam pwm_g_1_cry_9_c_inv_LC_2_30_1.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_9_c_inv_LC_2_30_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 pwm_g_1_cry_9_c_inv_LC_2_30_1 (
            .in0(_gnd_net_),
            .in1(N__3327),
            .in2(N__2525),
            .in3(N__2512),
            .lcout(pwm_ctr_i_9),
            .ltout(),
            .carryin(pwm_g_1_cry_8),
            .carryout(pwm_g_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_10_c_inv_LC_2_30_2.C_ON=1'b1;
    defparam pwm_g_1_cry_10_c_inv_LC_2_30_2.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_10_c_inv_LC_2_30_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 pwm_g_1_cry_10_c_inv_LC_2_30_2 (
            .in0(N__2500),
            .in1(N__3288),
            .in2(N__2666),
            .in3(_gnd_net_),
            .lcout(pwm_ctr_i_10),
            .ltout(),
            .carryin(pwm_g_1_cry_9),
            .carryout(pwm_g_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_1_cry_11_c_inv_LC_2_30_3.C_ON=1'b1;
    defparam pwm_g_1_cry_11_c_inv_LC_2_30_3.SEQ_MODE=4'b0000;
    defparam pwm_g_1_cry_11_c_inv_LC_2_30_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 pwm_g_1_cry_11_c_inv_LC_2_30_3 (
            .in0(N__2488),
            .in1(N__3252),
            .in2(N__2693),
            .in3(_gnd_net_),
            .lcout(pwm_ctr_i_11),
            .ltout(),
            .carryin(pwm_g_1_cry_10),
            .carryout(pwm_g_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_g_LC_2_30_4.C_ON=1'b0;
    defparam pwm_g_LC_2_30_4.SEQ_MODE=4'b1000;
    defparam pwm_g_LC_2_30_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_g_LC_2_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2681),
            .lcout(pwm_gZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3218),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_8_c_RNO_0_LC_2_30_5.C_ON=1'b0;
    defparam pwm_b_1_cry_8_c_RNO_0_LC_2_30_5.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_8_c_RNO_0_LC_2_30_5.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_8_c_RNO_0_LC_2_30_5 (
            .in0(N__4144),
            .in1(N__3803),
            .in2(_gnd_net_),
            .in3(N__3893),
            .lcout(),
            .ltout(N_71_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_8_c_RNO_LC_2_30_6.C_ON=1'b0;
    defparam pwm_b_1_cry_8_c_RNO_LC_2_30_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_8_c_RNO_LC_2_30_6.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_8_c_RNO_LC_2_30_6 (
            .in0(N__4423),
            .in1(N__3730),
            .in2(N__2669),
            .in3(N__4145),
            .lcout(pwm_b_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIKFG11_28_LC_2_30_7.C_ON=1'b0;
    defparam ctr_RNIKFG11_28_LC_2_30_7.SEQ_MODE=4'b0000;
    defparam ctr_RNIKFG11_28_LC_2_30_7.LUT_INIT=16'b0000010110100000;
    LogicCell40 ctr_RNIKFG11_28_LC_2_30_7 (
            .in0(N__3731),
            .in1(_gnd_net_),
            .in2(N__4224),
            .in3(N__4424),
            .lcout(pwm_g_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_0_c_LC_3_25_0.C_ON=1'b1;
    defparam un33_r_val_cry_0_c_LC_3_25_0.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_0_c_LC_3_25_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un33_r_val_cry_0_c_LC_3_25_0 (
            .in0(_gnd_net_),
            .in1(N__4865),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(un33_r_val_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_0_THRU_LUT4_0_LC_3_25_1.C_ON=1'b1;
    defparam un33_r_val_cry_0_THRU_LUT4_0_LC_3_25_1.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_0_THRU_LUT4_0_LC_3_25_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_0_THRU_LUT4_0_LC_3_25_1 (
            .in0(_gnd_net_),
            .in1(N__2656),
            .in2(N__2773),
            .in3(N__2639),
            .lcout(un33_r_val_cry_0_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_0),
            .carryout(un33_r_val_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_1_THRU_LUT4_0_LC_3_25_2.C_ON=1'b1;
    defparam un33_r_val_cry_1_THRU_LUT4_0_LC_3_25_2.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_1_THRU_LUT4_0_LC_3_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_1_THRU_LUT4_0_LC_3_25_2 (
            .in0(_gnd_net_),
            .in1(N__2755),
            .in2(N__4899),
            .in3(N__2636),
            .lcout(un33_r_val_cry_1_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_1),
            .carryout(un33_r_val_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_2_THRU_LUT4_0_LC_3_25_3.C_ON=1'b1;
    defparam un33_r_val_cry_2_THRU_LUT4_0_LC_3_25_3.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_2_THRU_LUT4_0_LC_3_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_2_THRU_LUT4_0_LC_3_25_3 (
            .in0(_gnd_net_),
            .in1(N__2758),
            .in2(N__3556),
            .in3(N__2633),
            .lcout(un33_r_val_cry_2_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_2),
            .carryout(un33_r_val_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_3_THRU_LUT4_0_LC_3_25_4.C_ON=1'b1;
    defparam un33_r_val_cry_3_THRU_LUT4_0_LC_3_25_4.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_3_THRU_LUT4_0_LC_3_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_3_THRU_LUT4_0_LC_3_25_4 (
            .in0(_gnd_net_),
            .in1(N__2756),
            .in2(N__3652),
            .in3(N__2822),
            .lcout(un33_r_val_cry_3_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_3),
            .carryout(un33_r_val_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_4_THRU_LUT4_0_LC_3_25_5.C_ON=1'b1;
    defparam un33_r_val_cry_4_THRU_LUT4_0_LC_3_25_5.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_4_THRU_LUT4_0_LC_3_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_4_THRU_LUT4_0_LC_3_25_5 (
            .in0(_gnd_net_),
            .in1(N__2759),
            .in2(N__3424),
            .in3(N__2810),
            .lcout(un33_r_val_cry_4_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_4),
            .carryout(un33_r_val_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_5_THRU_LUT4_0_LC_3_25_6.C_ON=1'b1;
    defparam un33_r_val_cry_5_THRU_LUT4_0_LC_3_25_6.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_5_THRU_LUT4_0_LC_3_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_5_THRU_LUT4_0_LC_3_25_6 (
            .in0(_gnd_net_),
            .in1(N__2757),
            .in2(N__3840),
            .in3(N__2807),
            .lcout(un33_r_val_cry_5_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_5),
            .carryout(un33_r_val_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_6_THRU_LUT4_0_LC_3_25_7.C_ON=1'b1;
    defparam un33_r_val_cry_6_THRU_LUT4_0_LC_3_25_7.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_6_THRU_LUT4_0_LC_3_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_6_THRU_LUT4_0_LC_3_25_7 (
            .in0(_gnd_net_),
            .in1(N__2760),
            .in2(N__4629),
            .in3(N__2804),
            .lcout(un33_r_val_cry_6_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_6),
            .carryout(un33_r_val_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_7_THRU_LUT4_0_LC_3_26_0.C_ON=1'b1;
    defparam un33_r_val_cry_7_THRU_LUT4_0_LC_3_26_0.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_7_THRU_LUT4_0_LC_3_26_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_7_THRU_LUT4_0_LC_3_26_0 (
            .in0(_gnd_net_),
            .in1(N__2761),
            .in2(N__3882),
            .in3(N__2801),
            .lcout(un33_r_val_cry_7_THRU_CO),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(un33_r_val_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_8_THRU_LUT4_0_LC_3_26_1.C_ON=1'b1;
    defparam un33_r_val_cry_8_THRU_LUT4_0_LC_3_26_1.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_8_THRU_LUT4_0_LC_3_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_8_THRU_LUT4_0_LC_3_26_1 (
            .in0(_gnd_net_),
            .in1(N__2762),
            .in2(N__3190),
            .in3(N__2711),
            .lcout(un33_r_val_cry_8_THRU_CO),
            .ltout(),
            .carryin(un33_r_val_cry_8),
            .carryout(un33_r_val_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_10_c_RNO_0_LC_3_26_2.C_ON=1'b1;
    defparam pwm_r_1_cry_10_c_RNO_0_LC_3_26_2.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_10_c_RNO_0_LC_3_26_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 pwm_r_1_cry_10_c_RNO_0_LC_3_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2879),
            .in3(N__2708),
            .lcout(pwm_r_1_cry_10_c_RNOZ0Z_0),
            .ltout(),
            .carryin(un33_r_val_cry_9),
            .carryout(un33_r_val_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un33_r_val_cry_10_THRU_LUT4_0_LC_3_26_3.C_ON=1'b0;
    defparam un33_r_val_cry_10_THRU_LUT4_0_LC_3_26_3.SEQ_MODE=4'b0000;
    defparam un33_r_val_cry_10_THRU_LUT4_0_LC_3_26_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un33_r_val_cry_10_THRU_LUT4_0_LC_3_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2705),
            .lcout(),
            .ltout(un33_r_val_cry_10_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_11_c_RNO_0_LC_3_26_4.C_ON=1'b0;
    defparam pwm_r_1_cry_11_c_RNO_0_LC_3_26_4.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_11_c_RNO_0_LC_3_26_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 pwm_r_1_cry_11_c_RNO_0_LC_3_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2702),
            .in3(N__2699),
            .lcout(pwm_r_1_cry_11_c_RNOZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_4_c_RNO_0_LC_3_26_5.C_ON=1'b0;
    defparam pwm_r_1_cry_4_c_RNO_0_LC_3_26_5.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_4_c_RNO_0_LC_3_26_5.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_4_c_RNO_0_LC_3_26_5 (
            .in0(N__4793),
            .in1(N__3648),
            .in2(N__4258),
            .in3(N__2864),
            .lcout(),
            .ltout(N_91_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_4_c_RNO_LC_3_26_6.C_ON=1'b0;
    defparam pwm_r_1_cry_4_c_RNO_LC_3_26_6.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_4_c_RNO_LC_3_26_6.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_4_c_RNO_LC_3_26_6 (
            .in0(N__4458),
            .in1(N__4221),
            .in2(N__2858),
            .in3(N__4726),
            .lcout(pwm_r_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_0_c_LC_3_27_0.C_ON=1'b1;
    defparam pwm_r_1_cry_0_c_LC_3_27_0.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_0_c_LC_3_27_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_0_c_LC_3_27_0 (
            .in0(_gnd_net_),
            .in1(N__2855),
            .in2(N__3149),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_27_0_),
            .carryout(pwm_r_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_1_c_LC_3_27_1.C_ON=1'b1;
    defparam pwm_r_1_cry_1_c_LC_3_27_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_1_c_LC_3_27_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_1_c_LC_3_27_1 (
            .in0(_gnd_net_),
            .in1(N__2849),
            .in2(N__3122),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_0),
            .carryout(pwm_r_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_2_c_LC_3_27_2.C_ON=1'b1;
    defparam pwm_r_1_cry_2_c_LC_3_27_2.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_2_c_LC_3_27_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_2_c_LC_3_27_2 (
            .in0(_gnd_net_),
            .in1(N__3083),
            .in2(N__3626),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_1),
            .carryout(pwm_r_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_3_c_LC_3_27_3.C_ON=1'b1;
    defparam pwm_r_1_cry_3_c_LC_3_27_3.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_3_c_LC_3_27_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_3_c_LC_3_27_3 (
            .in0(_gnd_net_),
            .in1(N__3050),
            .in2(N__3524),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_2),
            .carryout(pwm_r_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_4_c_LC_3_27_4.C_ON=1'b1;
    defparam pwm_r_1_cry_4_c_LC_3_27_4.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_4_c_LC_3_27_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_4_c_LC_3_27_4 (
            .in0(_gnd_net_),
            .in1(N__3026),
            .in2(N__2840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_3),
            .carryout(pwm_r_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_5_c_LC_3_27_5.C_ON=1'b1;
    defparam pwm_r_1_cry_5_c_LC_3_27_5.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_5_c_LC_3_27_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_5_c_LC_3_27_5 (
            .in0(_gnd_net_),
            .in1(N__2999),
            .in2(N__2831),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_4),
            .carryout(pwm_r_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_6_c_LC_3_27_6.C_ON=1'b1;
    defparam pwm_r_1_cry_6_c_LC_3_27_6.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_6_c_LC_3_27_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_6_c_LC_3_27_6 (
            .in0(_gnd_net_),
            .in1(N__2975),
            .in2(N__3503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_5),
            .carryout(pwm_r_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_7_c_LC_3_27_7.C_ON=1'b1;
    defparam pwm_r_1_cry_7_c_LC_3_27_7.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_7_c_LC_3_27_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_7_c_LC_3_27_7 (
            .in0(_gnd_net_),
            .in1(N__2945),
            .in2(N__3374),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_6),
            .carryout(pwm_r_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_8_c_LC_3_28_0.C_ON=1'b1;
    defparam pwm_r_1_cry_8_c_LC_3_28_0.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_8_c_LC_3_28_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_8_c_LC_3_28_0 (
            .in0(_gnd_net_),
            .in1(N__3359),
            .in2(N__3854),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_28_0_),
            .carryout(pwm_r_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_9_c_LC_3_28_1.C_ON=1'b1;
    defparam pwm_r_1_cry_9_c_LC_3_28_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_9_c_LC_3_28_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_9_c_LC_3_28_1 (
            .in0(_gnd_net_),
            .in1(N__3335),
            .in2(N__2888),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_8),
            .carryout(pwm_r_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_10_c_LC_3_28_2.C_ON=1'b1;
    defparam pwm_r_1_cry_10_c_LC_3_28_2.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_10_c_LC_3_28_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_10_c_LC_3_28_2 (
            .in0(_gnd_net_),
            .in1(N__3662),
            .in2(N__3302),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_9),
            .carryout(pwm_r_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_11_c_LC_3_28_3.C_ON=1'b1;
    defparam pwm_r_1_cry_11_c_LC_3_28_3.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_11_c_LC_3_28_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_r_1_cry_11_c_LC_3_28_3 (
            .in0(_gnd_net_),
            .in1(N__3262),
            .in2(N__3914),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_r_1_cry_10),
            .carryout(pwm_r_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_LC_3_28_4.C_ON=1'b0;
    defparam pwm_r_LC_3_28_4.SEQ_MODE=4'b1000;
    defparam pwm_r_LC_3_28_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_r_LC_3_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2915),
            .lcout(pwm_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3223),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_9_c_RNO_0_LC_3_28_5.C_ON=1'b0;
    defparam pwm_r_1_cry_9_c_RNO_0_LC_3_28_5.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_9_c_RNO_0_LC_3_28_5.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_9_c_RNO_0_LC_3_28_5 (
            .in0(N__4528),
            .in1(N__3186),
            .in2(N__4226),
            .in3(N__2900),
            .lcout(),
            .ltout(N_96_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_9_c_RNO_LC_3_28_6.C_ON=1'b0;
    defparam pwm_r_1_cry_9_c_RNO_LC_3_28_6.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_9_c_RNO_LC_3_28_6.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_9_c_RNO_LC_3_28_6 (
            .in0(N__4419),
            .in1(N__4159),
            .in2(N__2891),
            .in3(N__3981),
            .lcout(pwm_r_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_10_c_RNO_LC_3_28_7.C_ON=1'b0;
    defparam pwm_b_1_cry_10_c_RNO_LC_3_28_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_10_c_RNO_LC_3_28_7.LUT_INIT=16'b0000100011001000;
    LogicCell40 pwm_b_1_cry_10_c_RNO_LC_3_28_7 (
            .in0(N__3724),
            .in1(N__4418),
            .in2(N__4225),
            .in3(N__2878),
            .lcout(pwm_b_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_0_c_LC_3_29_0.C_ON=1'b1;
    defparam pwm_b_1_cry_0_c_LC_3_29_0.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_0_c_LC_3_29_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_0_c_LC_3_29_0 (
            .in0(_gnd_net_),
            .in1(N__4913),
            .in2(N__3148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(pwm_b_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_1_c_LC_3_29_1.C_ON=1'b1;
    defparam pwm_b_1_cry_1_c_LC_3_29_1.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_1_c_LC_3_29_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_1_c_LC_3_29_1 (
            .in0(_gnd_net_),
            .in1(N__3111),
            .in2(N__3092),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_0),
            .carryout(pwm_b_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_2_c_LC_3_29_2.C_ON=1'b1;
    defparam pwm_b_1_cry_2_c_LC_3_29_2.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_2_c_LC_3_29_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_2_c_LC_3_29_2 (
            .in0(_gnd_net_),
            .in1(N__4802),
            .in2(N__3082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_1),
            .carryout(pwm_b_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_3_c_LC_3_29_3.C_ON=1'b1;
    defparam pwm_b_1_cry_3_c_LC_3_29_3.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_3_c_LC_3_29_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_3_c_LC_3_29_3 (
            .in0(_gnd_net_),
            .in1(N__3059),
            .in2(N__3049),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_2),
            .carryout(pwm_b_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_4_c_LC_3_29_4.C_ON=1'b1;
    defparam pwm_b_1_cry_4_c_LC_3_29_4.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_4_c_LC_3_29_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_4_c_LC_3_29_4 (
            .in0(_gnd_net_),
            .in1(N__4949),
            .in2(N__3022),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_3),
            .carryout(pwm_b_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_5_c_LC_3_29_5.C_ON=1'b1;
    defparam pwm_b_1_cry_5_c_LC_3_29_5.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_5_c_LC_3_29_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_5_c_LC_3_29_5 (
            .in0(_gnd_net_),
            .in1(N__3398),
            .in2(N__2998),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_4),
            .carryout(pwm_b_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_6_c_LC_3_29_6.C_ON=1'b1;
    defparam pwm_b_1_cry_6_c_LC_3_29_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_6_c_LC_3_29_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_6_c_LC_3_29_6 (
            .in0(_gnd_net_),
            .in1(N__3746),
            .in2(N__2974),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_5),
            .carryout(pwm_b_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_7_c_LC_3_29_7.C_ON=1'b1;
    defparam pwm_b_1_cry_7_c_LC_3_29_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_7_c_LC_3_29_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_7_c_LC_3_29_7 (
            .in0(_gnd_net_),
            .in1(N__3992),
            .in2(N__2944),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_6),
            .carryout(pwm_b_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_8_c_LC_3_30_0.C_ON=1'b1;
    defparam pwm_b_1_cry_8_c_LC_3_30_0.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_8_c_LC_3_30_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_8_c_LC_3_30_0 (
            .in0(_gnd_net_),
            .in1(N__3365),
            .in2(N__3358),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_30_0_),
            .carryout(pwm_b_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_9_c_LC_3_30_1.C_ON=1'b1;
    defparam pwm_b_1_cry_9_c_LC_3_30_1.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_9_c_LC_3_30_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_9_c_LC_3_30_1 (
            .in0(_gnd_net_),
            .in1(N__3164),
            .in2(N__3334),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_8),
            .carryout(pwm_b_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_10_c_LC_3_30_2.C_ON=1'b1;
    defparam pwm_b_1_cry_10_c_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_10_c_LC_3_30_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_10_c_LC_3_30_2 (
            .in0(_gnd_net_),
            .in1(N__3311),
            .in2(N__3301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_9),
            .carryout(pwm_b_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_11_c_LC_3_30_3.C_ON=1'b1;
    defparam pwm_b_1_cry_11_c_LC_3_30_3.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_11_c_LC_3_30_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 pwm_b_1_cry_11_c_LC_3_30_3 (
            .in0(_gnd_net_),
            .in1(N__3272),
            .in2(N__3263),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(pwm_b_1_cry_10),
            .carryout(pwm_b_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_LC_3_30_4.C_ON=1'b0;
    defparam pwm_b_LC_3_30_4.SEQ_MODE=4'b1000;
    defparam pwm_b_LC_3_30_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_b_LC_3_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3236),
            .lcout(pwm_bZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3220),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_9_c_RNO_0_LC_3_30_6.C_ON=1'b0;
    defparam pwm_b_1_cry_9_c_RNO_0_LC_3_30_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_9_c_RNO_0_LC_3_30_6.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_9_c_RNO_0_LC_3_30_6 (
            .in0(N__4222),
            .in1(N__4539),
            .in2(_gnd_net_),
            .in3(N__3194),
            .lcout(),
            .ltout(N_72_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_9_c_RNO_LC_3_30_7.C_ON=1'b0;
    defparam pwm_b_1_cry_9_c_RNO_LC_3_30_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_9_c_RNO_LC_3_30_7.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_9_c_RNO_LC_3_30_7 (
            .in0(N__4459),
            .in1(N__4223),
            .in2(N__3167),
            .in3(N__3985),
            .lcout(pwm_b_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_2_c_RNO_0_LC_4_25_0.C_ON=1'b0;
    defparam pwm_r_1_cry_2_c_RNO_0_LC_4_25_0.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_2_c_RNO_0_LC_4_25_0.LUT_INIT=16'b0010111000011101;
    LogicCell40 pwm_r_1_cry_2_c_RNO_0_LC_4_25_0 (
            .in0(N__4906),
            .in1(N__4205),
            .in2(N__4873),
            .in3(N__3158),
            .lcout(),
            .ltout(N_89_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_2_c_RNO_LC_4_25_1.C_ON=1'b0;
    defparam pwm_r_1_cry_2_c_RNO_LC_4_25_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_2_c_RNO_LC_4_25_1.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_2_c_RNO_LC_4_25_1 (
            .in0(N__4434),
            .in1(N__4217),
            .in2(N__3152),
            .in3(N__4796),
            .lcout(pwm_r_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_3_c_RNO_0_LC_4_25_3.C_ON=1'b0;
    defparam pwm_r_1_cry_3_c_RNO_0_LC_4_25_3.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_3_c_RNO_0_LC_4_25_3.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_3_c_RNO_0_LC_4_25_3 (
            .in0(N__3613),
            .in1(N__3560),
            .in2(N__4254),
            .in3(N__3533),
            .lcout(),
            .ltout(N_90_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_3_c_RNO_LC_4_25_4.C_ON=1'b0;
    defparam pwm_r_1_cry_3_c_RNO_LC_4_25_4.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_3_c_RNO_LC_4_25_4.LUT_INIT=16'b1011100000110000;
    LogicCell40 pwm_r_1_cry_3_c_RNO_LC_4_25_4 (
            .in0(N__3494),
            .in1(N__4435),
            .in2(N__3527),
            .in3(N__4209),
            .lcout(pwm_r_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_6_c_RNO_0_LC_4_26_0.C_ON=1'b0;
    defparam pwm_r_1_cry_6_c_RNO_0_LC_4_26_0.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_6_c_RNO_0_LC_4_26_0.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_6_c_RNO_0_LC_4_26_0 (
            .in0(N__4724),
            .in1(N__3841),
            .in2(N__4259),
            .in3(N__3512),
            .lcout(),
            .ltout(N_93_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_6_c_RNO_LC_4_26_1.C_ON=1'b0;
    defparam pwm_r_1_cry_6_c_RNO_LC_4_26_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_6_c_RNO_LC_4_26_1.LUT_INIT=16'b1000100011110000;
    LogicCell40 pwm_r_1_cry_6_c_RNO_LC_4_26_1 (
            .in0(N__3812),
            .in1(N__4233),
            .in2(N__3506),
            .in3(N__4461),
            .lcout(pwm_r_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_5_c_RNO_0_LC_4_26_4.C_ON=1'b0;
    defparam pwm_b_1_cry_5_c_RNO_0_LC_4_26_4.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_5_c_RNO_0_LC_4_26_4.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_5_c_RNO_0_LC_4_26_4 (
            .in0(N__4227),
            .in1(N__3489),
            .in2(_gnd_net_),
            .in3(N__3425),
            .lcout(),
            .ltout(N_68_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_5_c_RNO_LC_4_26_5.C_ON=1'b0;
    defparam pwm_b_1_cry_5_c_RNO_LC_4_26_5.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_5_c_RNO_LC_4_26_5.LUT_INIT=16'b1100000011010001;
    LogicCell40 pwm_b_1_cry_5_c_RNO_LC_4_26_5 (
            .in0(N__4603),
            .in1(N__4460),
            .in2(N__3401),
            .in3(N__4228),
            .lcout(pwm_b_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_7_c_RNO_0_LC_4_26_6.C_ON=1'b0;
    defparam pwm_r_1_cry_7_c_RNO_0_LC_4_26_6.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_7_c_RNO_0_LC_4_26_6.LUT_INIT=16'b0111001000100111;
    LogicCell40 pwm_r_1_cry_7_c_RNO_0_LC_4_26_6 (
            .in0(N__4232),
            .in1(N__4604),
            .in2(N__3386),
            .in3(N__4633),
            .lcout(),
            .ltout(N_94_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_7_c_RNO_LC_4_26_7.C_ON=1'b0;
    defparam pwm_r_1_cry_7_c_RNO_LC_4_26_7.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_7_c_RNO_LC_4_26_7.LUT_INIT=16'b1000100011110000;
    LogicCell40 pwm_r_1_cry_7_c_RNO_LC_4_26_7 (
            .in0(N__4541),
            .in1(N__4234),
            .in2(N__3377),
            .in3(N__4462),
            .lcout(pwm_r_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_11_c_RNO_LC_4_27_1.C_ON=1'b0;
    defparam pwm_r_1_cry_11_c_RNO_LC_4_27_1.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_11_c_RNO_LC_4_27_1.LUT_INIT=16'b0001001100000010;
    LogicCell40 pwm_r_1_cry_11_c_RNO_LC_4_27_1 (
            .in0(N__4253),
            .in1(N__4442),
            .in2(N__3986),
            .in3(N__3920),
            .lcout(pwm_r_1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIP7LC1_24_LC_4_27_2.C_ON=1'b0;
    defparam ctr_RNIP7LC1_24_LC_4_27_2.SEQ_MODE=4'b0000;
    defparam ctr_RNIP7LC1_24_LC_4_27_2.LUT_INIT=16'b1101100000011011;
    LogicCell40 ctr_RNIP7LC1_24_LC_4_27_2 (
            .in0(N__4723),
            .in1(N__4244),
            .in2(N__4463),
            .in3(N__3805),
            .lcout(pwm_g_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_8_c_RNO_0_LC_4_27_3.C_ON=1'b0;
    defparam pwm_r_1_cry_8_c_RNO_0_LC_4_27_3.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_8_c_RNO_0_LC_4_27_3.LUT_INIT=16'b0101110001010011;
    LogicCell40 pwm_r_1_cry_8_c_RNO_0_LC_4_27_3 (
            .in0(N__3807),
            .in1(N__3889),
            .in2(N__4261),
            .in3(N__3863),
            .lcout(),
            .ltout(N_95_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_8_c_RNO_LC_4_27_4.C_ON=1'b0;
    defparam pwm_r_1_cry_8_c_RNO_LC_4_27_4.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_8_c_RNO_LC_4_27_4.LUT_INIT=16'b1101100001010000;
    LogicCell40 pwm_r_1_cry_8_c_RNO_LC_4_27_4 (
            .in0(N__4440),
            .in1(N__4249),
            .in2(N__3857),
            .in3(N__3735),
            .lcout(pwm_r_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_6_c_RNO_0_LC_4_27_5.C_ON=1'b0;
    defparam pwm_b_1_cry_6_c_RNO_0_LC_4_27_5.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_6_c_RNO_0_LC_4_27_5.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_6_c_RNO_0_LC_4_27_5 (
            .in0(N__4243),
            .in1(N__4722),
            .in2(_gnd_net_),
            .in3(N__3845),
            .lcout(),
            .ltout(N_69_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_6_c_RNO_LC_4_27_6.C_ON=1'b0;
    defparam pwm_b_1_cry_6_c_RNO_LC_4_27_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_6_c_RNO_LC_4_27_6.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_6_c_RNO_LC_4_27_6 (
            .in0(N__4439),
            .in1(N__4245),
            .in2(N__3815),
            .in3(N__3806),
            .lcout(pwm_b_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_r_1_cry_10_c_RNO_LC_4_27_7.C_ON=1'b0;
    defparam pwm_r_1_cry_10_c_RNO_LC_4_27_7.SEQ_MODE=4'b0000;
    defparam pwm_r_1_cry_10_c_RNO_LC_4_27_7.LUT_INIT=16'b0001001100010000;
    LogicCell40 pwm_r_1_cry_10_c_RNO_LC_4_27_7 (
            .in0(N__3736),
            .in1(N__4441),
            .in2(N__4262),
            .in3(N__3668),
            .lcout(pwm_r_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_4_c_RNO_0_LC_4_28_0.C_ON=1'b0;
    defparam pwm_b_1_cry_4_c_RNO_0_LC_4_28_0.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_4_c_RNO_0_LC_4_28_0.LUT_INIT=16'b0100010011101110;
    LogicCell40 pwm_b_1_cry_4_c_RNO_0_LC_4_28_0 (
            .in0(N__4255),
            .in1(N__4784),
            .in2(_gnd_net_),
            .in3(N__3656),
            .lcout(),
            .ltout(N_67_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_4_c_RNO_LC_4_28_1.C_ON=1'b0;
    defparam pwm_b_1_cry_4_c_RNO_LC_4_28_1.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_4_c_RNO_LC_4_28_1.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_4_c_RNO_LC_4_28_1 (
            .in0(N__4465),
            .in1(N__4257),
            .in2(N__3629),
            .in3(N__4725),
            .lcout(pwm_b_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_0_c_RNO_LC_4_28_7.C_ON=1'b0;
    defparam pwm_b_1_cry_0_c_RNO_LC_4_28_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_0_c_RNO_LC_4_28_7.LUT_INIT=16'b0000101010001101;
    LogicCell40 pwm_b_1_cry_0_c_RNO_LC_4_28_7 (
            .in0(N__4464),
            .in1(N__4943),
            .in2(N__4877),
            .in3(N__4256),
            .lcout(pwm_b_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_2_c_RNO_0_LC_4_29_0.C_ON=1'b0;
    defparam pwm_b_1_cry_2_c_RNO_0_LC_4_29_0.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_2_c_RNO_0_LC_4_29_0.LUT_INIT=16'b0111011100100010;
    LogicCell40 pwm_b_1_cry_2_c_RNO_0_LC_4_29_0 (
            .in0(N__4235),
            .in1(N__4907),
            .in2(_gnd_net_),
            .in3(N__4872),
            .lcout(),
            .ltout(N_65_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_2_c_RNO_LC_4_29_1.C_ON=1'b0;
    defparam pwm_b_1_cry_2_c_RNO_LC_4_29_1.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_2_c_RNO_LC_4_29_1.LUT_INIT=16'b1010000010110001;
    LogicCell40 pwm_b_1_cry_2_c_RNO_LC_4_29_1 (
            .in0(N__4471),
            .in1(N__4239),
            .in2(N__4805),
            .in3(N__4794),
            .lcout(pwm_b_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIL3LC1_22_LC_4_29_2.C_ON=1'b0;
    defparam ctr_RNIL3LC1_22_LC_4_29_2.SEQ_MODE=4'b0000;
    defparam ctr_RNIL3LC1_22_LC_4_29_2.LUT_INIT=16'b1110010000100111;
    LogicCell40 ctr_RNIL3LC1_22_LC_4_29_2 (
            .in0(N__4795),
            .in1(N__4470),
            .in2(N__4260),
            .in3(N__4727),
            .lcout(pwm_g_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ctr_RNIR9LC1_25_LC_4_29_4.C_ON=1'b0;
    defparam ctr_RNIR9LC1_25_LC_4_29_4.SEQ_MODE=4'b0000;
    defparam ctr_RNIR9LC1_25_LC_4_29_4.LUT_INIT=16'b1000101111010001;
    LogicCell40 ctr_RNIR9LC1_25_LC_4_29_4 (
            .in0(N__4240),
            .in1(N__4534),
            .in2(N__4472),
            .in3(N__4602),
            .lcout(pwm_g_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_7_c_RNO_0_LC_4_29_6.C_ON=1'b0;
    defparam pwm_b_1_cry_7_c_RNO_0_LC_4_29_6.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_7_c_RNO_0_LC_4_29_6.LUT_INIT=16'b0111011100100010;
    LogicCell40 pwm_b_1_cry_7_c_RNO_0_LC_4_29_6 (
            .in0(N__4241),
            .in1(N__4634),
            .in2(_gnd_net_),
            .in3(N__4601),
            .lcout(),
            .ltout(N_70_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_b_1_cry_7_c_RNO_LC_4_29_7.C_ON=1'b0;
    defparam pwm_b_1_cry_7_c_RNO_LC_4_29_7.SEQ_MODE=4'b0000;
    defparam pwm_b_1_cry_7_c_RNO_LC_4_29_7.LUT_INIT=16'b1100000011010001;
    LogicCell40 pwm_b_1_cry_7_c_RNO_LC_4_29_7 (
            .in0(N__4535),
            .in1(N__4469),
            .in2(N__4265),
            .in3(N__4242),
            .lcout(pwm_b_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
